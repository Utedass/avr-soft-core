<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-55.2452,20.0193,101.958,-57.6833</PageViewport>
<gate>
<ID>1</ID>
<type>DA_FROM</type>
<position>-26,-12.5</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID R16_LD</lparam></gate>
<gate>
<ID>2</ID>
<type>DA_FROM</type>
<position>-26,-18.5</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID R16_ALU_A</lparam></gate>
<gate>
<ID>3</ID>
<type>DA_FROM</type>
<position>-26,-21.5</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID R16_ALU_B</lparam></gate>
<gate>
<ID>4</ID>
<type>DA_FROM</type>
<position>-26,-15.5</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID R16_DATA</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>-30,-12.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>-30,-15.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_TOGGLE</type>
<position>-30,-18.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>-30,-21.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>9</ID>
<type>DA_FROM</type>
<position>-26,-26.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID R17_LD</lparam></gate>
<gate>
<ID>10</ID>
<type>DA_FROM</type>
<position>-26,-32.5</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID R17_ALU_A</lparam></gate>
<gate>
<ID>11</ID>
<type>DA_FROM</type>
<position>-26,-35.5</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID R17_ALU_B</lparam></gate>
<gate>
<ID>12</ID>
<type>DA_FROM</type>
<position>-26,-29.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID R17_DATA</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>-30,-26.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>-30,-29.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>-30,-32.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>-30,-35.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>17</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>-31.5,15.5</position>
<input>
<ID>ENABLE_0</ID>10 </input>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>20 </input>
<input>
<ID>IN_2</ID>21 </input>
<input>
<ID>IN_3</ID>22 </input>
<input>
<ID>IN_4</ID>23 </input>
<input>
<ID>IN_5</ID>24 </input>
<input>
<ID>IN_6</ID>25 </input>
<input>
<ID>IN_7</ID>26 </input>
<output>
<ID>OUT_0</ID>11 </output>
<output>
<ID>OUT_1</ID>12 </output>
<output>
<ID>OUT_2</ID>13 </output>
<output>
<ID>OUT_3</ID>18 </output>
<output>
<ID>OUT_4</ID>14 </output>
<output>
<ID>OUT_5</ID>17 </output>
<output>
<ID>OUT_6</ID>15 </output>
<output>
<ID>OUT_7</ID>16 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>18</ID>
<type>DA_FROM</type>
<position>-38.5,15.5</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MANUAL_DATA</lparam></gate>
<gate>
<ID>19</ID>
<type>DE_TO</type>
<position>-28,19.5</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>20</ID>
<type>DE_TO</type>
<position>-29,24.5</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>21</ID>
<type>DE_TO</type>
<position>-30,19.5</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>22</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>73,-101</position>
<output>
<ID>A_equal_B</ID>33 </output>
<output>
<ID>A_greater_B</ID>32 </output>
<output>
<ID>A_less_B</ID>34 </output>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>68 </input>
<input>
<ID>IN_2</ID>69 </input>
<input>
<ID>IN_3</ID>70 </input>
<input>
<ID>IN_B_0</ID>51 </input>
<input>
<ID>IN_B_1</ID>52 </input>
<input>
<ID>IN_B_2</ID>53 </input>
<input>
<ID>IN_B_3</ID>54 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>23</ID>
<type>DE_TO</type>
<position>-32,19.5</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_FULLADDER_4BIT</type>
<position>92,-100.5</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_2</ID>73 </input>
<input>
<ID>IN_3</ID>74 </input>
<input>
<ID>IN_B_0</ID>55 </input>
<input>
<ID>IN_B_1</ID>56 </input>
<input>
<ID>IN_B_2</ID>57 </input>
<input>
<ID>IN_B_3</ID>58 </input>
<input>
<ID>carry_in</ID>9 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>25</ID>
<type>AE_FULLADDER_4BIT</type>
<position>108,-100.5</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>68 </input>
<input>
<ID>IN_2</ID>69 </input>
<input>
<ID>IN_3</ID>70 </input>
<input>
<ID>IN_B_0</ID>51 </input>
<input>
<ID>IN_B_1</ID>52 </input>
<input>
<ID>IN_B_2</ID>53 </input>
<input>
<ID>IN_B_3</ID>54 </input>
<output>
<ID>carry_out</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>26</ID>
<type>DE_TO</type>
<position>-34,19.5</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>27</ID>
<type>DE_TO</type>
<position>-31,24.5</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>28</ID>
<type>DE_TO</type>
<position>-33,24.5</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>29</ID>
<type>DE_TO</type>
<position>-35,24.5</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>31</ID>
<type>DD_KEYPAD_HEX</type>
<position>-65.5,8</position>
<output>
<ID>OUT_0</ID>23 </output>
<output>
<ID>OUT_1</ID>24 </output>
<output>
<ID>OUT_2</ID>25 </output>
<output>
<ID>OUT_3</ID>26 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>32</ID>
<type>DD_KEYPAD_HEX</type>
<position>-53.5,8</position>
<output>
<ID>OUT_0</ID>19 </output>
<output>
<ID>OUT_1</ID>20 </output>
<output>
<ID>OUT_2</ID>21 </output>
<output>
<ID>OUT_3</ID>22 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>33</ID>
<type>DA_FROM</type>
<position>-26,-7.5</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID MANUAL_DATA</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>-30,-7.5</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>43</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>57,-101</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_2</ID>73 </input>
<input>
<ID>IN_3</ID>74 </input>
<input>
<ID>IN_B_0</ID>55 </input>
<input>
<ID>IN_B_1</ID>56 </input>
<input>
<ID>IN_B_2</ID>57 </input>
<input>
<ID>IN_B_3</ID>58 </input>
<input>
<ID>in_A_equal_B</ID>33 </input>
<input>
<ID>in_A_greater_B</ID>32 </input>
<input>
<ID>in_A_less_B</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>47</ID>
<type>HA_JUNC_2</type>
<position>78,-81</position>
<input>
<ID>N_in1</ID>58 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>48</ID>
<type>HA_JUNC_2</type>
<position>79,-81</position>
<input>
<ID>N_in1</ID>57 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>49</ID>
<type>HA_JUNC_2</type>
<position>80,-81</position>
<input>
<ID>N_in1</ID>56 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>50</ID>
<type>HA_JUNC_2</type>
<position>81,-81</position>
<input>
<ID>N_in1</ID>55 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>51</ID>
<type>HA_JUNC_2</type>
<position>82,-81</position>
<input>
<ID>N_in1</ID>54 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>52</ID>
<type>AE_REGISTER8</type>
<position>30,5</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>65 </input>
<input>
<ID>IN_2</ID>59 </input>
<input>
<ID>IN_3</ID>63 </input>
<input>
<ID>IN_4</ID>62 </input>
<input>
<ID>IN_5</ID>60 </input>
<input>
<ID>IN_6</ID>64 </input>
<input>
<ID>IN_7</ID>66 </input>
<output>
<ID>OUT_0</ID>80 </output>
<output>
<ID>OUT_1</ID>81 </output>
<output>
<ID>OUT_2</ID>82 </output>
<output>
<ID>OUT_3</ID>83 </output>
<output>
<ID>OUT_4</ID>84 </output>
<output>
<ID>OUT_5</ID>85 </output>
<output>
<ID>OUT_6</ID>86 </output>
<output>
<ID>OUT_7</ID>87 </output>
<input>
<ID>clear</ID>77 </input>
<input>
<ID>clock</ID>156 </input>
<input>
<ID>load</ID>76 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 18</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>53</ID>
<type>HA_JUNC_2</type>
<position>83,-81</position>
<input>
<ID>N_in1</ID>53 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>54</ID>
<type>HA_JUNC_2</type>
<position>7,90.5</position>
<input>
<ID>N_in0</ID>120 </input>
<input>
<ID>N_in1</ID>66 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>55</ID>
<type>HA_JUNC_2</type>
<position>8,90.5</position>
<input>
<ID>N_in0</ID>116 </input>
<input>
<ID>N_in1</ID>64 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>56</ID>
<type>HA_JUNC_2</type>
<position>9,90.5</position>
<input>
<ID>N_in0</ID>119 </input>
<input>
<ID>N_in1</ID>60 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>57</ID>
<type>HA_JUNC_2</type>
<position>10,90.5</position>
<input>
<ID>N_in0</ID>115 </input>
<input>
<ID>N_in1</ID>62 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>58</ID>
<type>HA_JUNC_2</type>
<position>11,90.5</position>
<input>
<ID>N_in0</ID>118 </input>
<input>
<ID>N_in1</ID>63 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>59</ID>
<type>HA_JUNC_2</type>
<position>12,90.5</position>
<input>
<ID>N_in0</ID>113 </input>
<input>
<ID>N_in1</ID>59 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>60</ID>
<type>HA_JUNC_2</type>
<position>13,90.5</position>
<input>
<ID>N_in0</ID>117 </input>
<input>
<ID>N_in1</ID>65 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>61</ID>
<type>HA_JUNC_2</type>
<position>14,90.5</position>
<input>
<ID>N_in0</ID>114 </input>
<input>
<ID>N_in1</ID>61 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>62</ID>
<type>HA_JUNC_2</type>
<position>7,-121</position>
<input>
<ID>N_in0</ID>66 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>63</ID>
<type>HA_JUNC_2</type>
<position>8,-121</position>
<input>
<ID>N_in0</ID>64 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>64</ID>
<type>HA_JUNC_2</type>
<position>9,-121</position>
<input>
<ID>N_in0</ID>60 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>65</ID>
<type>HA_JUNC_2</type>
<position>10,-121</position>
<input>
<ID>N_in0</ID>62 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>66</ID>
<type>HA_JUNC_2</type>
<position>11,-121</position>
<input>
<ID>N_in0</ID>63 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>67</ID>
<type>HA_JUNC_2</type>
<position>12,-121</position>
<input>
<ID>N_in0</ID>59 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>68</ID>
<type>HA_JUNC_2</type>
<position>13,-121</position>
<input>
<ID>N_in0</ID>65 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>69</ID>
<type>HA_JUNC_2</type>
<position>14,-121</position>
<input>
<ID>N_in0</ID>61 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>70</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>86.5,12</position>
<input>
<ID>ENABLE_0</ID>79 </input>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>81 </input>
<input>
<ID>IN_2</ID>82 </input>
<input>
<ID>IN_3</ID>83 </input>
<input>
<ID>IN_4</ID>84 </input>
<input>
<ID>IN_5</ID>85 </input>
<input>
<ID>IN_6</ID>86 </input>
<input>
<ID>IN_7</ID>87 </input>
<output>
<ID>OUT_0</ID>99 </output>
<output>
<ID>OUT_1</ID>103 </output>
<output>
<ID>OUT_2</ID>100 </output>
<output>
<ID>OUT_3</ID>104 </output>
<output>
<ID>OUT_4</ID>101 </output>
<output>
<ID>OUT_5</ID>108 </output>
<output>
<ID>OUT_6</ID>102 </output>
<output>
<ID>OUT_7</ID>107 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>71</ID>
<type>HA_JUNC_2</type>
<position>84,-81</position>
<input>
<ID>N_in1</ID>52 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>72</ID>
<type>HA_JUNC_2</type>
<position>85,-81</position>
<input>
<ID>N_in1</ID>51 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>73</ID>
<type>HA_JUNC_2</type>
<position>66,-81</position>
<input>
<ID>N_in1</ID>74 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>30.5,17.5</position>
<gparam>LABEL_TEXT R16</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>HA_JUNC_2</type>
<position>67,-81</position>
<input>
<ID>N_in1</ID>73 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>76</ID>
<type>DA_FROM</type>
<position>26.5,12.5</position>
<input>
<ID>IN_0</ID>76 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R16_LD</lparam></gate>
<gate>
<ID>77</ID>
<type>DA_FROM</type>
<position>29,-3.5</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R16_CLR</lparam></gate>
<gate>
<ID>78</ID>
<type>DA_FROM</type>
<position>79.5,12</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R16_ALU_A</lparam></gate>
<gate>
<ID>79</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>110.5,12</position>
<input>
<ID>ENABLE_0</ID>88 </input>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>81 </input>
<input>
<ID>IN_2</ID>82 </input>
<input>
<ID>IN_3</ID>83 </input>
<input>
<ID>IN_4</ID>84 </input>
<input>
<ID>IN_5</ID>85 </input>
<input>
<ID>IN_6</ID>86 </input>
<input>
<ID>IN_7</ID>87 </input>
<output>
<ID>OUT_0</ID>110 </output>
<output>
<ID>OUT_2</ID>109 </output>
<output>
<ID>OUT_4</ID>111 </output>
<output>
<ID>OUT_6</ID>112 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>80</ID>
<type>DA_FROM</type>
<position>103.5,12</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R16_ALU_B</lparam></gate>
<gate>
<ID>81</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>62,12</position>
<input>
<ID>ENABLE_0</ID>89 </input>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>81 </input>
<input>
<ID>IN_2</ID>82 </input>
<input>
<ID>IN_3</ID>83 </input>
<input>
<ID>IN_4</ID>84 </input>
<input>
<ID>IN_5</ID>85 </input>
<input>
<ID>IN_6</ID>86 </input>
<input>
<ID>IN_7</ID>87 </input>
<output>
<ID>OUT_0</ID>90 </output>
<output>
<ID>OUT_1</ID>91 </output>
<output>
<ID>OUT_2</ID>92 </output>
<output>
<ID>OUT_3</ID>98 </output>
<output>
<ID>OUT_4</ID>93 </output>
<output>
<ID>OUT_5</ID>97 </output>
<output>
<ID>OUT_6</ID>94 </output>
<output>
<ID>OUT_7</ID>96 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>82</ID>
<type>DA_FROM</type>
<position>55,12</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R16_DATA</lparam></gate>
<gate>
<ID>83</ID>
<type>HA_JUNC_2</type>
<position>68,-81</position>
<input>
<ID>N_in1</ID>72 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>84</ID>
<type>HA_JUNC_2</type>
<position>69,-81</position>
<input>
<ID>N_in1</ID>71 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>85</ID>
<type>DE_TO</type>
<position>65.5,16</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>86</ID>
<type>DE_TO</type>
<position>64.5,21</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>87</ID>
<type>DE_TO</type>
<position>63.5,16</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>88</ID>
<type>DE_TO</type>
<position>61.5,16</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>89</ID>
<type>DE_TO</type>
<position>59.5,16</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>90</ID>
<type>HA_JUNC_2</type>
<position>70,-81</position>
<input>
<ID>N_in1</ID>70 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>91</ID>
<type>DE_TO</type>
<position>62.5,21</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>92</ID>
<type>DE_TO</type>
<position>60.5,21</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>93</ID>
<type>DE_TO</type>
<position>58.5,21</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>94</ID>
<type>DE_TO</type>
<position>90,16</position>
<input>
<ID>IN_0</ID>99 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A0</lparam></gate>
<gate>
<ID>95</ID>
<type>DE_TO</type>
<position>88,16</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A2</lparam></gate>
<gate>
<ID>96</ID>
<type>DE_TO</type>
<position>86,16</position>
<input>
<ID>IN_0</ID>101 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A4</lparam></gate>
<gate>
<ID>97</ID>
<type>DE_TO</type>
<position>84,16</position>
<input>
<ID>IN_0</ID>102 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A6</lparam></gate>
<gate>
<ID>98</ID>
<type>DE_TO</type>
<position>89,26.5</position>
<input>
<ID>IN_0</ID>103 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A1</lparam></gate>
<gate>
<ID>99</ID>
<type>DE_TO</type>
<position>87,26.5</position>
<input>
<ID>IN_0</ID>104 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A3</lparam></gate>
<gate>
<ID>100</ID>
<type>DE_TO</type>
<position>85,26.5</position>
<input>
<ID>IN_0</ID>108 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A5</lparam></gate>
<gate>
<ID>101</ID>
<type>DE_TO</type>
<position>83,26.5</position>
<input>
<ID>IN_0</ID>107 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A7</lparam></gate>
<gate>
<ID>102</ID>
<type>DE_TO</type>
<position>114,16</position>
<input>
<ID>IN_0</ID>110 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B0</lparam></gate>
<gate>
<ID>103</ID>
<type>DE_TO</type>
<position>112,16</position>
<input>
<ID>IN_0</ID>109 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B2</lparam></gate>
<gate>
<ID>104</ID>
<type>DE_TO</type>
<position>110,16</position>
<input>
<ID>IN_0</ID>111 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B4</lparam></gate>
<gate>
<ID>105</ID>
<type>DE_TO</type>
<position>108,16</position>
<input>
<ID>IN_0</ID>112 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B6</lparam></gate>
<gate>
<ID>106</ID>
<type>DE_TO</type>
<position>113,26.5</position>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B1</lparam></gate>
<gate>
<ID>107</ID>
<type>DE_TO</type>
<position>111,26.5</position>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B3</lparam></gate>
<gate>
<ID>108</ID>
<type>DE_TO</type>
<position>109,26.5</position>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B5</lparam></gate>
<gate>
<ID>109</ID>
<type>DE_TO</type>
<position>107,26.5</position>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B7</lparam></gate>
<gate>
<ID>110</ID>
<type>DE_TO</type>
<position>14,93.5</position>
<input>
<ID>IN_0</ID>114 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>111</ID>
<type>DE_TO</type>
<position>13,98.5</position>
<input>
<ID>IN_0</ID>117 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>112</ID>
<type>DE_TO</type>
<position>12,93.5</position>
<input>
<ID>IN_0</ID>113 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>113</ID>
<type>DE_TO</type>
<position>10,93.5</position>
<input>
<ID>IN_0</ID>115 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>114</ID>
<type>DE_TO</type>
<position>8,93.5</position>
<input>
<ID>IN_0</ID>116 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>115</ID>
<type>DE_TO</type>
<position>11,98.5</position>
<input>
<ID>IN_0</ID>118 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>116</ID>
<type>DE_TO</type>
<position>9,98.5</position>
<input>
<ID>IN_0</ID>119 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>117</ID>
<type>DE_TO</type>
<position>7,98.5</position>
<input>
<ID>IN_0</ID>120 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>118</ID>
<type>HA_JUNC_2</type>
<position>71,-81</position>
<input>
<ID>N_in1</ID>69 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>119</ID>
<type>HA_JUNC_2</type>
<position>72,-81</position>
<input>
<ID>N_in1</ID>68 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>120</ID>
<type>HA_JUNC_2</type>
<position>73,-81</position>
<input>
<ID>N_in1</ID>67 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>121</ID>
<type>AE_REGISTER8</type>
<position>30,-33.5</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>65 </input>
<input>
<ID>IN_2</ID>59 </input>
<input>
<ID>IN_3</ID>63 </input>
<input>
<ID>IN_4</ID>62 </input>
<input>
<ID>IN_5</ID>60 </input>
<input>
<ID>IN_6</ID>64 </input>
<input>
<ID>IN_7</ID>66 </input>
<output>
<ID>OUT_0</ID>125 </output>
<output>
<ID>OUT_1</ID>126 </output>
<output>
<ID>OUT_2</ID>127 </output>
<output>
<ID>OUT_3</ID>128 </output>
<output>
<ID>OUT_4</ID>129 </output>
<output>
<ID>OUT_5</ID>130 </output>
<output>
<ID>OUT_6</ID>131 </output>
<output>
<ID>OUT_7</ID>132 </output>
<input>
<ID>clear</ID>123 </input>
<input>
<ID>clock</ID>155 </input>
<input>
<ID>load</ID>122 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>122</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>86.5,-26.5</position>
<input>
<ID>ENABLE_0</ID>124 </input>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>126 </input>
<input>
<ID>IN_2</ID>127 </input>
<input>
<ID>IN_3</ID>128 </input>
<input>
<ID>IN_4</ID>129 </input>
<input>
<ID>IN_5</ID>130 </input>
<input>
<ID>IN_6</ID>131 </input>
<input>
<ID>IN_7</ID>132 </input>
<output>
<ID>OUT_0</ID>143 </output>
<output>
<ID>OUT_1</ID>147 </output>
<output>
<ID>OUT_2</ID>144 </output>
<output>
<ID>OUT_3</ID>148 </output>
<output>
<ID>OUT_4</ID>145 </output>
<output>
<ID>OUT_5</ID>150 </output>
<output>
<ID>OUT_6</ID>146 </output>
<output>
<ID>OUT_7</ID>149 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_LABEL</type>
<position>30.5,-21</position>
<gparam>LABEL_TEXT R17</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>124</ID>
<type>DA_FROM</type>
<position>26.5,-26</position>
<input>
<ID>IN_0</ID>122 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R17_LD</lparam></gate>
<gate>
<ID>125</ID>
<type>DA_FROM</type>
<position>29,-41.5</position>
<input>
<ID>IN_0</ID>123 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R17_CLR</lparam></gate>
<gate>
<ID>126</ID>
<type>DA_FROM</type>
<position>79.5,-26.5</position>
<input>
<ID>IN_0</ID>124 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R17_ALU_A</lparam></gate>
<gate>
<ID>127</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>110.5,-26.5</position>
<input>
<ID>ENABLE_0</ID>133 </input>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>126 </input>
<input>
<ID>IN_2</ID>127 </input>
<input>
<ID>IN_3</ID>128 </input>
<input>
<ID>IN_4</ID>129 </input>
<input>
<ID>IN_5</ID>130 </input>
<input>
<ID>IN_6</ID>131 </input>
<input>
<ID>IN_7</ID>132 </input>
<output>
<ID>OUT_0</ID>152 </output>
<output>
<ID>OUT_2</ID>151 </output>
<output>
<ID>OUT_4</ID>153 </output>
<output>
<ID>OUT_6</ID>154 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>128</ID>
<type>DA_FROM</type>
<position>103.5,-26.5</position>
<input>
<ID>IN_0</ID>133 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R17_ALU_B</lparam></gate>
<gate>
<ID>129</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>62,-26.5</position>
<input>
<ID>ENABLE_0</ID>134 </input>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>126 </input>
<input>
<ID>IN_2</ID>127 </input>
<input>
<ID>IN_3</ID>128 </input>
<input>
<ID>IN_4</ID>129 </input>
<input>
<ID>IN_5</ID>130 </input>
<input>
<ID>IN_6</ID>131 </input>
<input>
<ID>IN_7</ID>132 </input>
<output>
<ID>OUT_0</ID>135 </output>
<output>
<ID>OUT_1</ID>136 </output>
<output>
<ID>OUT_2</ID>137 </output>
<output>
<ID>OUT_3</ID>142 </output>
<output>
<ID>OUT_4</ID>138 </output>
<output>
<ID>OUT_5</ID>141 </output>
<output>
<ID>OUT_6</ID>139 </output>
<output>
<ID>OUT_7</ID>140 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>130</ID>
<type>DA_FROM</type>
<position>55,-26.5</position>
<input>
<ID>IN_0</ID>134 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R17_DATA</lparam></gate>
<gate>
<ID>131</ID>
<type>DE_TO</type>
<position>65.5,-22.5</position>
<input>
<ID>IN_0</ID>135 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>132</ID>
<type>DE_TO</type>
<position>64.5,-17.5</position>
<input>
<ID>IN_0</ID>136 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>133</ID>
<type>DE_TO</type>
<position>63.5,-22.5</position>
<input>
<ID>IN_0</ID>137 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>134</ID>
<type>DE_TO</type>
<position>61.5,-22.5</position>
<input>
<ID>IN_0</ID>138 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>135</ID>
<type>DE_TO</type>
<position>59.5,-22.5</position>
<input>
<ID>IN_0</ID>139 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>136</ID>
<type>DE_TO</type>
<position>62.5,-17.5</position>
<input>
<ID>IN_0</ID>142 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>137</ID>
<type>DE_TO</type>
<position>60.5,-17.5</position>
<input>
<ID>IN_0</ID>141 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>138</ID>
<type>DE_TO</type>
<position>58.5,-17.5</position>
<input>
<ID>IN_0</ID>140 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>139</ID>
<type>DE_TO</type>
<position>90,-22.5</position>
<input>
<ID>IN_0</ID>143 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A0</lparam></gate>
<gate>
<ID>140</ID>
<type>DE_TO</type>
<position>88,-22.5</position>
<input>
<ID>IN_0</ID>144 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A2</lparam></gate>
<gate>
<ID>141</ID>
<type>DE_TO</type>
<position>86,-22.5</position>
<input>
<ID>IN_0</ID>145 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A4</lparam></gate>
<gate>
<ID>142</ID>
<type>DE_TO</type>
<position>84,-22.5</position>
<input>
<ID>IN_0</ID>146 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A6</lparam></gate>
<gate>
<ID>143</ID>
<type>DE_TO</type>
<position>89,-12</position>
<input>
<ID>IN_0</ID>147 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A1</lparam></gate>
<gate>
<ID>144</ID>
<type>DE_TO</type>
<position>87,-12</position>
<input>
<ID>IN_0</ID>148 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A3</lparam></gate>
<gate>
<ID>145</ID>
<type>DE_TO</type>
<position>85,-12</position>
<input>
<ID>IN_0</ID>150 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A5</lparam></gate>
<gate>
<ID>146</ID>
<type>DE_TO</type>
<position>83,-12</position>
<input>
<ID>IN_0</ID>149 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A7</lparam></gate>
<gate>
<ID>147</ID>
<type>DE_TO</type>
<position>114,-22.5</position>
<input>
<ID>IN_0</ID>152 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B0</lparam></gate>
<gate>
<ID>148</ID>
<type>DE_TO</type>
<position>112,-22.5</position>
<input>
<ID>IN_0</ID>151 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B2</lparam></gate>
<gate>
<ID>149</ID>
<type>DE_TO</type>
<position>110,-22.5</position>
<input>
<ID>IN_0</ID>153 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B4</lparam></gate>
<gate>
<ID>150</ID>
<type>DE_TO</type>
<position>108,-22.5</position>
<input>
<ID>IN_0</ID>154 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B6</lparam></gate>
<gate>
<ID>151</ID>
<type>DE_TO</type>
<position>113,-12</position>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B1</lparam></gate>
<gate>
<ID>152</ID>
<type>DE_TO</type>
<position>111,-12</position>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B3</lparam></gate>
<gate>
<ID>153</ID>
<type>DE_TO</type>
<position>109,-12</position>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B5</lparam></gate>
<gate>
<ID>154</ID>
<type>DE_TO</type>
<position>107,-12</position>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B7</lparam></gate>
<gate>
<ID>155</ID>
<type>DA_FROM</type>
<position>27,-39.5</position>
<input>
<ID>IN_0</ID>155 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>156</ID>
<type>DA_FROM</type>
<position>27,-1</position>
<input>
<ID>IN_0</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>157</ID>
<type>DA_FROM</type>
<position>-26,-3</position>
<input>
<ID>IN_0</ID>157 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_TOGGLE</type>
<position>-30,-3</position>
<output>
<ID>OUT_0</ID>157 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-12.5,-28,-12.5</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-28,-12.5,-28,-12.5</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>-28 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-15.5,-28,-15.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-18.5,-28,-18.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-28,-18.5,-28,-18.5</points>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection>
<intersection>-28 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-21.5,-28,-21.5</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-26.5,-28,-26.5</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-29.5,-28,-29.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-32.5,-28,-32.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-35.5,-28,-35.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>100,-99.5,100,-99.5</points>
<connection>
<GID>24</GID>
<name>carry_in</name></connection>
<connection>
<GID>25</GID>
<name>carry_out</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,15.5,-36.5,15.5</points>
<connection>
<GID>17</GID>
<name>ENABLE_0</name></connection>
<intersection>15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-36.5,15.5,-36.5,15.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,17.5,-28,17.5</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<connection>
<GID>19</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,17.5,-29,22.5</points>
<connection>
<GID>17</GID>
<name>OUT_1</name></connection>
<connection>
<GID>20</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,17.5,-30,17.5</points>
<connection>
<GID>17</GID>
<name>OUT_2</name></connection>
<connection>
<GID>21</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32,17.5,-32,17.5</points>
<connection>
<GID>17</GID>
<name>OUT_4</name></connection>
<connection>
<GID>23</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,17.5,-34,17.5</points>
<connection>
<GID>17</GID>
<name>OUT_6</name></connection>
<connection>
<GID>26</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,17.5,-35,22.5</points>
<connection>
<GID>17</GID>
<name>OUT_7</name></connection>
<connection>
<GID>29</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33,17.5,-33,22.5</points>
<connection>
<GID>17</GID>
<name>OUT_5</name></connection>
<connection>
<GID>28</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31,17.5,-31,22.5</points>
<connection>
<GID>17</GID>
<name>OUT_3</name></connection>
<connection>
<GID>27</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,5,-28,13.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48.5,5,-28,5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>-28 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,7,-29,13.5</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48.5,7,-29,7</points>
<connection>
<GID>32</GID>
<name>OUT_1</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,9,-30,13.5</points>
<connection>
<GID>17</GID>
<name>IN_2</name></connection>
<intersection>9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48.5,9,-30,9</points>
<connection>
<GID>32</GID>
<name>OUT_2</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31,11,-31,13.5</points>
<connection>
<GID>17</GID>
<name>IN_3</name></connection>
<intersection>11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48.5,11,-31,11</points>
<connection>
<GID>32</GID>
<name>OUT_3</name></connection>
<intersection>-31 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32,0,-32,13.5</points>
<connection>
<GID>17</GID>
<name>IN_4</name></connection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-60,0,-32,0</points>
<intersection>-60 2</intersection>
<intersection>-32 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-60,0,-60,5</points>
<intersection>0 1</intersection>
<intersection>5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-60.5,5,-60,5</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>-60 2</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33,0.5,-33,13.5</points>
<connection>
<GID>17</GID>
<name>IN_5</name></connection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-59.5,0.5,-33,0.5</points>
<intersection>-59.5 2</intersection>
<intersection>-33 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-59.5,0.5,-59.5,7</points>
<intersection>0.5 1</intersection>
<intersection>7 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-60.5,7,-59.5,7</points>
<connection>
<GID>31</GID>
<name>OUT_1</name></connection>
<intersection>-59.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,1,-34,13.5</points>
<connection>
<GID>17</GID>
<name>IN_6</name></connection>
<intersection>1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-59,1,-34,1</points>
<intersection>-59 2</intersection>
<intersection>-34 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-59,1,-59,9</points>
<intersection>1 1</intersection>
<intersection>9 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-60.5,9,-59,9</points>
<connection>
<GID>31</GID>
<name>OUT_2</name></connection>
<intersection>-59 2</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,1.5,-35,13.5</points>
<connection>
<GID>17</GID>
<name>IN_7</name></connection>
<intersection>1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-58.5,1.5,-35,1.5</points>
<intersection>-58.5 2</intersection>
<intersection>-35 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-58.5,1.5,-58.5,11</points>
<intersection>1.5 1</intersection>
<intersection>11 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-60.5,11,-58.5,11</points>
<connection>
<GID>31</GID>
<name>OUT_3</name></connection>
<intersection>-58.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-7.5,-28,-7.5</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>65,-99,65,-99</points>
<connection>
<GID>22</GID>
<name>A_greater_B</name></connection>
<connection>
<GID>43</GID>
<name>in_A_greater_B</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>65,-101,65,-101</points>
<connection>
<GID>22</GID>
<name>A_equal_B</name></connection>
<connection>
<GID>43</GID>
<name>in_A_equal_B</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>65,-103,65,-103</points>
<connection>
<GID>22</GID>
<name>A_less_B</name></connection>
<connection>
<GID>43</GID>
<name>in_A_less_B</name></connection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,-96.5,113,-91.5</points>
<connection>
<GID>25</GID>
<name>IN_B_0</name></connection>
<intersection>-91.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>85,-91.5,85,-82</points>
<connection>
<GID>72</GID>
<name>N_in1</name></connection>
<intersection>-91.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>78,-91.5,113,-91.5</points>
<intersection>78 7</intersection>
<intersection>85 1</intersection>
<intersection>113 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>78,-97,78,-91.5</points>
<connection>
<GID>22</GID>
<name>IN_B_0</name></connection>
<intersection>-91.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-91,84,-82</points>
<connection>
<GID>71</GID>
<name>N_in1</name></connection>
<intersection>-91 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>112,-96.5,112,-91</points>
<connection>
<GID>25</GID>
<name>IN_B_1</name></connection>
<intersection>-91 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>77,-91,112,-91</points>
<intersection>77 7</intersection>
<intersection>84 0</intersection>
<intersection>112 1</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>77,-97,77,-91</points>
<connection>
<GID>22</GID>
<name>IN_B_1</name></connection>
<intersection>-91 2</intersection></vsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-96.5,111,-90.5</points>
<connection>
<GID>25</GID>
<name>IN_B_2</name></connection>
<intersection>-90.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>83,-90.5,83,-82</points>
<connection>
<GID>53</GID>
<name>N_in1</name></connection>
<intersection>-90.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>76,-90.5,111,-90.5</points>
<intersection>76 7</intersection>
<intersection>83 1</intersection>
<intersection>111 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>76,-97,76,-90.5</points>
<connection>
<GID>22</GID>
<name>IN_B_2</name></connection>
<intersection>-90.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-90,82,-82</points>
<connection>
<GID>51</GID>
<name>N_in1</name></connection>
<intersection>-90 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>110,-96.5,110,-90</points>
<connection>
<GID>25</GID>
<name>IN_B_3</name></connection>
<intersection>-90 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>75,-90,110,-90</points>
<intersection>75 7</intersection>
<intersection>82 0</intersection>
<intersection>110 1</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>75,-97,75,-90</points>
<connection>
<GID>22</GID>
<name>IN_B_3</name></connection>
<intersection>-90 2</intersection></vsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-96.5,97,-89.5</points>
<connection>
<GID>24</GID>
<name>IN_B_0</name></connection>
<intersection>-89.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>81,-89.5,81,-82</points>
<connection>
<GID>50</GID>
<name>N_in1</name></connection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>62,-89.5,97,-89.5</points>
<intersection>62 7</intersection>
<intersection>81 1</intersection>
<intersection>97 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>62,-97,62,-89.5</points>
<connection>
<GID>43</GID>
<name>IN_B_0</name></connection>
<intersection>-89.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-89,80,-82</points>
<connection>
<GID>49</GID>
<name>N_in1</name></connection>
<intersection>-89 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>96,-96.5,96,-89</points>
<connection>
<GID>24</GID>
<name>IN_B_1</name></connection>
<intersection>-89 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>61,-89,96,-89</points>
<intersection>61 7</intersection>
<intersection>80 0</intersection>
<intersection>96 1</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>61,-97,61,-89</points>
<connection>
<GID>43</GID>
<name>IN_B_1</name></connection>
<intersection>-89 2</intersection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95,-96.5,95,-88.5</points>
<connection>
<GID>24</GID>
<name>IN_B_2</name></connection>
<intersection>-88.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>79,-88.5,79,-82</points>
<connection>
<GID>48</GID>
<name>N_in1</name></connection>
<intersection>-88.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>60,-88.5,95,-88.5</points>
<intersection>60 7</intersection>
<intersection>79 1</intersection>
<intersection>95 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>60,-97,60,-88.5</points>
<connection>
<GID>43</GID>
<name>IN_B_2</name></connection>
<intersection>-88.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-88,78,-82</points>
<connection>
<GID>47</GID>
<name>N_in1</name></connection>
<intersection>-88 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>94,-96.5,94,-88</points>
<connection>
<GID>24</GID>
<name>IN_B_3</name></connection>
<intersection>-88 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>59,-88,94,-88</points>
<intersection>59 4</intersection>
<intersection>78 0</intersection>
<intersection>94 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>59,-97,59,-88</points>
<connection>
<GID>43</GID>
<name>IN_B_3</name></connection>
<intersection>-88 2</intersection></vsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-120,12,89.5</points>
<connection>
<GID>67</GID>
<name>N_in0</name></connection>
<connection>
<GID>59</GID>
<name>N_in1</name></connection>
<intersection>-34.5 8</intersection>
<intersection>4 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>12,4,26,4</points>
<connection>
<GID>52</GID>
<name>IN_2</name></connection>
<intersection>12 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>12,-34.5,26,-34.5</points>
<connection>
<GID>121</GID>
<name>IN_2</name></connection>
<intersection>12 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-120,9,89.5</points>
<connection>
<GID>64</GID>
<name>N_in0</name></connection>
<connection>
<GID>56</GID>
<name>N_in1</name></connection>
<intersection>-31.5 8</intersection>
<intersection>7 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>9,7,26,7</points>
<connection>
<GID>52</GID>
<name>IN_5</name></connection>
<intersection>9 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>9,-31.5,26,-31.5</points>
<connection>
<GID>121</GID>
<name>IN_5</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-120,14,89.5</points>
<connection>
<GID>69</GID>
<name>N_in0</name></connection>
<connection>
<GID>61</GID>
<name>N_in1</name></connection>
<intersection>-36.5 8</intersection>
<intersection>2 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>14,2,26,2</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>14,-36.5,26,-36.5</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-120,10,89.5</points>
<connection>
<GID>65</GID>
<name>N_in0</name></connection>
<connection>
<GID>57</GID>
<name>N_in1</name></connection>
<intersection>-32.5 8</intersection>
<intersection>6 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>10,6,26,6</points>
<connection>
<GID>52</GID>
<name>IN_4</name></connection>
<intersection>10 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>10,-32.5,26,-32.5</points>
<connection>
<GID>121</GID>
<name>IN_4</name></connection>
<intersection>10 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-120,11,89.5</points>
<connection>
<GID>66</GID>
<name>N_in0</name></connection>
<connection>
<GID>58</GID>
<name>N_in1</name></connection>
<intersection>-33.5 8</intersection>
<intersection>5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>11,5,26,5</points>
<connection>
<GID>52</GID>
<name>IN_3</name></connection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>11,-33.5,26,-33.5</points>
<connection>
<GID>121</GID>
<name>IN_3</name></connection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-120,8,89.5</points>
<connection>
<GID>63</GID>
<name>N_in0</name></connection>
<connection>
<GID>55</GID>
<name>N_in1</name></connection>
<intersection>-30.5 8</intersection>
<intersection>8 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>8,8,26,8</points>
<connection>
<GID>52</GID>
<name>IN_6</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>8,-30.5,26,-30.5</points>
<connection>
<GID>121</GID>
<name>IN_6</name></connection>
<intersection>8 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-120,13,89.5</points>
<connection>
<GID>68</GID>
<name>N_in0</name></connection>
<connection>
<GID>60</GID>
<name>N_in1</name></connection>
<intersection>-35.5 8</intersection>
<intersection>3 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>13,3,26,3</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>13,-35.5,26,-35.5</points>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<intersection>13 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-120,7,89.5</points>
<connection>
<GID>62</GID>
<name>N_in0</name></connection>
<connection>
<GID>54</GID>
<name>N_in1</name></connection>
<intersection>-29.5 8</intersection>
<intersection>9 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>7,9,26,9</points>
<connection>
<GID>52</GID>
<name>IN_7</name></connection>
<intersection>7 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>7,-29.5,26,-29.5</points>
<connection>
<GID>121</GID>
<name>IN_7</name></connection>
<intersection>7 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,-96.5,106,-86.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-86.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>73,-86.5,73,-82</points>
<connection>
<GID>120</GID>
<name>N_in1</name></connection>
<intersection>-86.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>71,-86.5,106,-86.5</points>
<intersection>71 4</intersection>
<intersection>73 1</intersection>
<intersection>106 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>71,-97,71,-86.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-86.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-86,72,-82</points>
<connection>
<GID>119</GID>
<name>N_in1</name></connection>
<intersection>-86 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>105,-96.5,105,-86</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>-86 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>70,-86,105,-86</points>
<intersection>70 4</intersection>
<intersection>72 0</intersection>
<intersection>105 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>70,-97,70,-86</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>-86 2</intersection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-96.5,104,-85.5</points>
<connection>
<GID>25</GID>
<name>IN_2</name></connection>
<intersection>-85.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>71,-85.5,71,-82</points>
<connection>
<GID>118</GID>
<name>N_in1</name></connection>
<intersection>-85.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>69,-85.5,104,-85.5</points>
<intersection>69 4</intersection>
<intersection>71 1</intersection>
<intersection>104 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>69,-97,69,-85.5</points>
<connection>
<GID>22</GID>
<name>IN_2</name></connection>
<intersection>-85.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-85,70,-82</points>
<connection>
<GID>90</GID>
<name>N_in1</name></connection>
<intersection>-85 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>103,-96.5,103,-85</points>
<connection>
<GID>25</GID>
<name>IN_3</name></connection>
<intersection>-85 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>68,-85,103,-85</points>
<intersection>68 4</intersection>
<intersection>70 0</intersection>
<intersection>103 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>68,-97,68,-85</points>
<connection>
<GID>22</GID>
<name>IN_3</name></connection>
<intersection>-85 2</intersection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-96.5,90,-84.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-84.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>69,-84.5,69,-82</points>
<connection>
<GID>84</GID>
<name>N_in1</name></connection>
<intersection>-84.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>55,-84.5,90,-84.5</points>
<intersection>55 4</intersection>
<intersection>69 1</intersection>
<intersection>90 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>55,-97,55,-84.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>-84.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-84,68,-82</points>
<connection>
<GID>83</GID>
<name>N_in1</name></connection>
<intersection>-84 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>89,-96.5,89,-84</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>-84 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>54,-84,89,-84</points>
<intersection>54 4</intersection>
<intersection>68 0</intersection>
<intersection>89 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>54,-97,54,-84</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>-84 2</intersection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-96.5,88,-83.5</points>
<connection>
<GID>24</GID>
<name>IN_2</name></connection>
<intersection>-83.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>67,-83.5,67,-82</points>
<connection>
<GID>75</GID>
<name>N_in1</name></connection>
<intersection>-83.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>53,-83.5,88,-83.5</points>
<intersection>53 4</intersection>
<intersection>67 1</intersection>
<intersection>88 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>53,-97,53,-83.5</points>
<connection>
<GID>43</GID>
<name>IN_2</name></connection>
<intersection>-83.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,-83,66,-82</points>
<connection>
<GID>73</GID>
<name>N_in1</name></connection>
<intersection>-83 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>87,-96.5,87,-83</points>
<connection>
<GID>24</GID>
<name>IN_3</name></connection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>52,-83,87,-83</points>
<intersection>52 4</intersection>
<intersection>66 0</intersection>
<intersection>87 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>52,-97,52,-83</points>
<connection>
<GID>43</GID>
<name>IN_3</name></connection>
<intersection>-83 2</intersection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,11,29,12.5</points>
<connection>
<GID>52</GID>
<name>load</name></connection>
<intersection>12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,12.5,29,12.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-3.5,31,0</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<connection>
<GID>52</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,12,81.5,12</points>
<connection>
<GID>70</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>78</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,2,90,10</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,2,114,2</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>65.5 4</intersection>
<intersection>90 0</intersection>
<intersection>114 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>114,2,114,10</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>2 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>65.5,2,65.5,10</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>2 1</intersection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,3,89,10</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>3 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,3,113,3</points>
<connection>
<GID>52</GID>
<name>OUT_1</name></connection>
<intersection>64.5 4</intersection>
<intersection>89 0</intersection>
<intersection>113 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>113,3,113,10</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>3 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>64.5,3,64.5,10</points>
<connection>
<GID>81</GID>
<name>IN_1</name></connection>
<intersection>3 1</intersection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,4,88,10</points>
<connection>
<GID>70</GID>
<name>IN_2</name></connection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,4,112,4</points>
<connection>
<GID>52</GID>
<name>OUT_2</name></connection>
<intersection>63.5 4</intersection>
<intersection>88 0</intersection>
<intersection>112 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>112,4,112,10</points>
<connection>
<GID>79</GID>
<name>IN_2</name></connection>
<intersection>4 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>63.5,4,63.5,10</points>
<connection>
<GID>81</GID>
<name>IN_2</name></connection>
<intersection>4 1</intersection></vsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,5,87,10</points>
<connection>
<GID>70</GID>
<name>IN_3</name></connection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,5,111,5</points>
<connection>
<GID>52</GID>
<name>OUT_3</name></connection>
<intersection>62.5 4</intersection>
<intersection>87 0</intersection>
<intersection>111 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>111,5,111,10</points>
<connection>
<GID>79</GID>
<name>IN_3</name></connection>
<intersection>5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>62.5,5,62.5,10</points>
<connection>
<GID>81</GID>
<name>IN_3</name></connection>
<intersection>5 1</intersection></vsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,6,86,10</points>
<connection>
<GID>70</GID>
<name>IN_4</name></connection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,6,110,6</points>
<connection>
<GID>52</GID>
<name>OUT_4</name></connection>
<intersection>61.5 4</intersection>
<intersection>86 0</intersection>
<intersection>110 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>110,6,110,10</points>
<connection>
<GID>79</GID>
<name>IN_4</name></connection>
<intersection>6 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>61.5,6,61.5,10</points>
<connection>
<GID>81</GID>
<name>IN_4</name></connection>
<intersection>6 1</intersection></vsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,7,85,10</points>
<connection>
<GID>70</GID>
<name>IN_5</name></connection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,7,109,7</points>
<connection>
<GID>52</GID>
<name>OUT_5</name></connection>
<intersection>60.5 4</intersection>
<intersection>85 0</intersection>
<intersection>109 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>109,7,109,10</points>
<connection>
<GID>79</GID>
<name>IN_5</name></connection>
<intersection>7 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>60.5,7,60.5,10</points>
<connection>
<GID>81</GID>
<name>IN_5</name></connection>
<intersection>7 1</intersection></vsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,8,84,10</points>
<connection>
<GID>70</GID>
<name>IN_6</name></connection>
<intersection>8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,8,108,8</points>
<connection>
<GID>52</GID>
<name>OUT_6</name></connection>
<intersection>59.5 5</intersection>
<intersection>84 0</intersection>
<intersection>108 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>108,8,108,10</points>
<connection>
<GID>79</GID>
<name>IN_6</name></connection>
<intersection>8 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>59.5,8,59.5,10</points>
<connection>
<GID>81</GID>
<name>IN_6</name></connection>
<intersection>8 1</intersection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,9,107,9</points>
<connection>
<GID>52</GID>
<name>OUT_7</name></connection>
<intersection>58.5 8</intersection>
<intersection>83 4</intersection>
<intersection>107 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>83,9,83,10</points>
<connection>
<GID>70</GID>
<name>IN_7</name></connection>
<intersection>9 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>107,9,107,10</points>
<connection>
<GID>79</GID>
<name>IN_7</name></connection>
<intersection>9 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>58.5,9,58.5,10</points>
<connection>
<GID>81</GID>
<name>IN_7</name></connection>
<intersection>9 1</intersection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,12,105.5,12</points>
<connection>
<GID>79</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>80</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,12,57,12</points>
<connection>
<GID>81</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>82</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,14,65.5,14</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<connection>
<GID>85</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,14,64.5,19</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<connection>
<GID>81</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,14,63.5,14</points>
<connection>
<GID>81</GID>
<name>OUT_2</name></connection>
<connection>
<GID>87</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,14,61.5,14</points>
<connection>
<GID>81</GID>
<name>OUT_4</name></connection>
<connection>
<GID>88</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,14,59.5,14</points>
<connection>
<GID>81</GID>
<name>OUT_6</name></connection>
<connection>
<GID>89</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,14,58.5,19</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<connection>
<GID>81</GID>
<name>OUT_7</name></connection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,14,60.5,19</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<connection>
<GID>81</GID>
<name>OUT_5</name></connection></vsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,14,62.5,19</points>
<connection>
<GID>81</GID>
<name>OUT_3</name></connection>
<connection>
<GID>91</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,14,90,14</points>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<connection>
<GID>94</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,14,88,14</points>
<connection>
<GID>70</GID>
<name>OUT_2</name></connection>
<connection>
<GID>95</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,14,86,14</points>
<connection>
<GID>70</GID>
<name>OUT_4</name></connection>
<connection>
<GID>96</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,14,84,14</points>
<connection>
<GID>70</GID>
<name>OUT_6</name></connection>
<connection>
<GID>97</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,14,89,24.5</points>
<connection>
<GID>70</GID>
<name>OUT_1</name></connection>
<connection>
<GID>98</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,14,87,24.5</points>
<connection>
<GID>70</GID>
<name>OUT_3</name></connection>
<connection>
<GID>99</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,14,83,24.5</points>
<connection>
<GID>70</GID>
<name>OUT_7</name></connection>
<connection>
<GID>101</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,14,85,24.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<connection>
<GID>70</GID>
<name>OUT_5</name></connection></vsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,14,112,14</points>
<connection>
<GID>79</GID>
<name>OUT_2</name></connection>
<connection>
<GID>103</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,14,114,14</points>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection>
<connection>
<GID>102</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,14,110,14</points>
<connection>
<GID>79</GID>
<name>OUT_4</name></connection>
<connection>
<GID>104</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,14,108,14</points>
<connection>
<GID>79</GID>
<name>OUT_6</name></connection>
<connection>
<GID>105</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,91.5,12,91.5</points>
<connection>
<GID>59</GID>
<name>N_in0</name></connection>
<connection>
<GID>112</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,91.5,14,91.5</points>
<connection>
<GID>61</GID>
<name>N_in0</name></connection>
<connection>
<GID>110</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,91.5,10,91.5</points>
<connection>
<GID>57</GID>
<name>N_in0</name></connection>
<connection>
<GID>113</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,91.5,8,91.5</points>
<connection>
<GID>55</GID>
<name>N_in0</name></connection>
<connection>
<GID>114</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,91.5,13,96.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<connection>
<GID>60</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,91.5,11,96.5</points>
<connection>
<GID>58</GID>
<name>N_in0</name></connection>
<connection>
<GID>115</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,91.5,9,96.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<connection>
<GID>56</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,91.5,7,96.5</points>
<connection>
<GID>54</GID>
<name>N_in0</name></connection>
<connection>
<GID>117</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-27.5,29,-26</points>
<connection>
<GID>121</GID>
<name>load</name></connection>
<intersection>-26 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>28.5,-26,29,-26</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-41.5,31,-38.5</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<connection>
<GID>121</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-26.5,81.5,-26.5</points>
<connection>
<GID>122</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>126</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-36.5,90,-28.5</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-36.5,114,-36.5</points>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection>
<intersection>65.5 4</intersection>
<intersection>90 0</intersection>
<intersection>114 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>114,-36.5,114,-28.5</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>-36.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>65.5,-36.5,65.5,-28.5</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<intersection>-36.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-35.5,89,-28.5</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-35.5,113,-35.5</points>
<connection>
<GID>121</GID>
<name>OUT_1</name></connection>
<intersection>64.5 4</intersection>
<intersection>89 0</intersection>
<intersection>113 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>113,-35.5,113,-28.5</points>
<connection>
<GID>127</GID>
<name>IN_1</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>64.5,-35.5,64.5,-28.5</points>
<connection>
<GID>129</GID>
<name>IN_1</name></connection>
<intersection>-35.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-34.5,88,-28.5</points>
<connection>
<GID>122</GID>
<name>IN_2</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-34.5,112,-34.5</points>
<connection>
<GID>121</GID>
<name>OUT_2</name></connection>
<intersection>63.5 4</intersection>
<intersection>88 0</intersection>
<intersection>112 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>112,-34.5,112,-28.5</points>
<connection>
<GID>127</GID>
<name>IN_2</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>63.5,-34.5,63.5,-28.5</points>
<connection>
<GID>129</GID>
<name>IN_2</name></connection>
<intersection>-34.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-33.5,87,-28.5</points>
<connection>
<GID>122</GID>
<name>IN_3</name></connection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-33.5,111,-33.5</points>
<connection>
<GID>121</GID>
<name>OUT_3</name></connection>
<intersection>62.5 4</intersection>
<intersection>87 0</intersection>
<intersection>111 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>111,-33.5,111,-28.5</points>
<connection>
<GID>127</GID>
<name>IN_3</name></connection>
<intersection>-33.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>62.5,-33.5,62.5,-28.5</points>
<connection>
<GID>129</GID>
<name>IN_3</name></connection>
<intersection>-33.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-32.5,86,-28.5</points>
<connection>
<GID>122</GID>
<name>IN_4</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-32.5,110,-32.5</points>
<connection>
<GID>121</GID>
<name>OUT_4</name></connection>
<intersection>61.5 4</intersection>
<intersection>86 0</intersection>
<intersection>110 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>110,-32.5,110,-28.5</points>
<connection>
<GID>127</GID>
<name>IN_4</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>61.5,-32.5,61.5,-28.5</points>
<connection>
<GID>129</GID>
<name>IN_4</name></connection>
<intersection>-32.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-31.5,85,-28.5</points>
<connection>
<GID>122</GID>
<name>IN_5</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-31.5,109,-31.5</points>
<connection>
<GID>121</GID>
<name>OUT_5</name></connection>
<intersection>60.5 4</intersection>
<intersection>85 0</intersection>
<intersection>109 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>109,-31.5,109,-28.5</points>
<connection>
<GID>127</GID>
<name>IN_5</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>60.5,-31.5,60.5,-28.5</points>
<connection>
<GID>129</GID>
<name>IN_5</name></connection>
<intersection>-31.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-30.5,84,-28.5</points>
<connection>
<GID>122</GID>
<name>IN_6</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-30.5,108,-30.5</points>
<connection>
<GID>121</GID>
<name>OUT_6</name></connection>
<intersection>59.5 5</intersection>
<intersection>84 0</intersection>
<intersection>108 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>108,-30.5,108,-28.5</points>
<connection>
<GID>127</GID>
<name>IN_6</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>59.5,-30.5,59.5,-28.5</points>
<connection>
<GID>129</GID>
<name>IN_6</name></connection>
<intersection>-30.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-29.5,107,-29.5</points>
<connection>
<GID>121</GID>
<name>OUT_7</name></connection>
<intersection>58.5 8</intersection>
<intersection>83 4</intersection>
<intersection>107 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>83,-29.5,83,-28.5</points>
<connection>
<GID>122</GID>
<name>IN_7</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>107,-29.5,107,-28.5</points>
<connection>
<GID>127</GID>
<name>IN_7</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>58.5,-29.5,58.5,-28.5</points>
<connection>
<GID>129</GID>
<name>IN_7</name></connection>
<intersection>-29.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-26.5,105.5,-26.5</points>
<connection>
<GID>127</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>128</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-26.5,57,-26.5</points>
<connection>
<GID>129</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>130</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-24.5,65.5,-24.5</points>
<connection>
<GID>129</GID>
<name>OUT_0</name></connection>
<connection>
<GID>131</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-24.5,64.5,-19.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<connection>
<GID>129</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-24.5,63.5,-24.5</points>
<connection>
<GID>129</GID>
<name>OUT_2</name></connection>
<connection>
<GID>133</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-24.5,61.5,-24.5</points>
<connection>
<GID>129</GID>
<name>OUT_4</name></connection>
<connection>
<GID>134</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-24.5,59.5,-24.5</points>
<connection>
<GID>129</GID>
<name>OUT_6</name></connection>
<connection>
<GID>135</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-24.5,58.5,-19.5</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<connection>
<GID>129</GID>
<name>OUT_7</name></connection></vsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-24.5,60.5,-19.5</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<connection>
<GID>129</GID>
<name>OUT_5</name></connection></vsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-24.5,62.5,-19.5</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<connection>
<GID>129</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-24.5,90,-24.5</points>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<connection>
<GID>139</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-24.5,88,-24.5</points>
<connection>
<GID>122</GID>
<name>OUT_2</name></connection>
<connection>
<GID>140</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-24.5,86,-24.5</points>
<connection>
<GID>122</GID>
<name>OUT_4</name></connection>
<connection>
<GID>141</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-24.5,84,-24.5</points>
<connection>
<GID>122</GID>
<name>OUT_6</name></connection>
<connection>
<GID>142</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-24.5,89,-14</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<connection>
<GID>122</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-24.5,87,-14</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<connection>
<GID>122</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-24.5,83,-14</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<connection>
<GID>122</GID>
<name>OUT_7</name></connection></vsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-24.5,85,-14</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<connection>
<GID>122</GID>
<name>OUT_5</name></connection></vsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-24.5,112,-24.5</points>
<connection>
<GID>127</GID>
<name>OUT_2</name></connection>
<connection>
<GID>148</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,-24.5,114,-24.5</points>
<connection>
<GID>127</GID>
<name>OUT_0</name></connection>
<connection>
<GID>147</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-24.5,110,-24.5</points>
<connection>
<GID>127</GID>
<name>OUT_4</name></connection>
<connection>
<GID>149</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-24.5,108,-24.5</points>
<connection>
<GID>127</GID>
<name>OUT_6</name></connection>
<connection>
<GID>150</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-39.5,29,-38.5</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<connection>
<GID>121</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-1,29,0</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<connection>
<GID>52</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-3,-28,-3</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<connection>
<GID>159</GID>
<name>OUT_0</name></connection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-8.42641e-006,1.25829,153.345,-74.537</PageViewport></page 1>
<page 2>
<PageViewport>-8.42641e-006,1.25829,153.345,-74.537</PageViewport></page 2>
<page 3>
<PageViewport>-8.42641e-006,1.25829,153.345,-74.537</PageViewport></page 3>
<page 4>
<PageViewport>-8.42641e-006,1.25829,153.345,-74.537</PageViewport></page 4>
<page 5>
<PageViewport>-8.42641e-006,1.25829,153.345,-74.537</PageViewport></page 5>
<page 6>
<PageViewport>-8.42641e-006,1.25829,153.345,-74.537</PageViewport></page 6>
<page 7>
<PageViewport>-8.42641e-006,1.25829,153.345,-74.537</PageViewport></page 7>
<page 8>
<PageViewport>-8.42641e-006,1.25829,153.345,-74.537</PageViewport></page 8>
<page 9>
<PageViewport>-8.42641e-006,1.25829,153.345,-74.537</PageViewport></page 9></circuit>
<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-53.5948,4.94504,284.973,-184.092</PageViewport>
<gate>
<ID>1</ID>
<type>DA_FROM</type>
<position>-26,-17</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID R16_LD</lparam></gate>
<gate>
<ID>4</ID>
<type>DA_FROM</type>
<position>-28,-104.5</position>
<input>
<ID>IN_0</ID>240 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID R16_DATA</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>-30,-17</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>9</ID>
<type>DA_FROM</type>
<position>-26,-20</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID R17_LD</lparam></gate>
<gate>
<ID>12</ID>
<type>DA_FROM</type>
<position>-14,-103.5</position>
<input>
<ID>IN_0</ID>236 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID R17_DATA</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>-30,-20</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>17</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>-31.5,15.5</position>
<input>
<ID>ENABLE_0</ID>10 </input>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>20 </input>
<input>
<ID>IN_2</ID>21 </input>
<input>
<ID>IN_3</ID>22 </input>
<input>
<ID>IN_4</ID>23 </input>
<input>
<ID>IN_5</ID>24 </input>
<input>
<ID>IN_6</ID>25 </input>
<input>
<ID>IN_7</ID>26 </input>
<output>
<ID>OUT_0</ID>11 </output>
<output>
<ID>OUT_1</ID>12 </output>
<output>
<ID>OUT_2</ID>13 </output>
<output>
<ID>OUT_3</ID>18 </output>
<output>
<ID>OUT_4</ID>14 </output>
<output>
<ID>OUT_5</ID>17 </output>
<output>
<ID>OUT_6</ID>15 </output>
<output>
<ID>OUT_7</ID>16 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>18</ID>
<type>DA_FROM</type>
<position>-38.5,15.5</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID MANUAL_DATA</lparam></gate>
<gate>
<ID>19</ID>
<type>DE_TO</type>
<position>-28,19.5</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>20</ID>
<type>DE_TO</type>
<position>-29,24.5</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>21</ID>
<type>DE_TO</type>
<position>-30,19.5</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>22</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>93,-100.5</position>
<output>
<ID>A_equal_B</ID>33 </output>
<output>
<ID>A_greater_B</ID>32 </output>
<output>
<ID>A_less_B</ID>34 </output>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>68 </input>
<input>
<ID>IN_2</ID>69 </input>
<input>
<ID>IN_3</ID>70 </input>
<input>
<ID>IN_B_0</ID>51 </input>
<input>
<ID>IN_B_1</ID>52 </input>
<input>
<ID>IN_B_2</ID>53 </input>
<input>
<ID>IN_B_3</ID>54 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>23</ID>
<type>DE_TO</type>
<position>-32,19.5</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>24</ID>
<type>AE_FULLADDER_4BIT</type>
<position>112,-100</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_2</ID>73 </input>
<input>
<ID>IN_3</ID>74 </input>
<input>
<ID>IN_B_0</ID>55 </input>
<input>
<ID>IN_B_1</ID>56 </input>
<input>
<ID>IN_B_2</ID>57 </input>
<input>
<ID>IN_B_3</ID>58 </input>
<output>
<ID>OUT_0</ID>167 </output>
<output>
<ID>OUT_1</ID>168 </output>
<output>
<ID>OUT_2</ID>169 </output>
<output>
<ID>OUT_3</ID>170 </output>
<input>
<ID>carry_in</ID>9 </input>
<output>
<ID>carry_out</ID>50 </output>
<output>
<ID>overflow</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>25</ID>
<type>AE_FULLADDER_4BIT</type>
<position>128,-100</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>68 </input>
<input>
<ID>IN_2</ID>69 </input>
<input>
<ID>IN_3</ID>70 </input>
<input>
<ID>IN_B_0</ID>51 </input>
<input>
<ID>IN_B_1</ID>52 </input>
<input>
<ID>IN_B_2</ID>53 </input>
<input>
<ID>IN_B_3</ID>54 </input>
<output>
<ID>OUT_0</ID>163 </output>
<output>
<ID>OUT_1</ID>164 </output>
<output>
<ID>OUT_2</ID>165 </output>
<output>
<ID>OUT_3</ID>166 </output>
<input>
<ID>carry_in</ID>75 </input>
<output>
<ID>carry_out</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>26</ID>
<type>DE_TO</type>
<position>-34,19.5</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>27</ID>
<type>DE_TO</type>
<position>-31,24.5</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>28</ID>
<type>DE_TO</type>
<position>-33,24.5</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>29</ID>
<type>DE_TO</type>
<position>-35,24.5</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>31</ID>
<type>DD_KEYPAD_HEX</type>
<position>-65.5,8</position>
<output>
<ID>OUT_0</ID>23 </output>
<output>
<ID>OUT_1</ID>24 </output>
<output>
<ID>OUT_2</ID>25 </output>
<output>
<ID>OUT_3</ID>26 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>32</ID>
<type>DD_KEYPAD_HEX</type>
<position>-53.5,8</position>
<output>
<ID>OUT_0</ID>19 </output>
<output>
<ID>OUT_1</ID>20 </output>
<output>
<ID>OUT_2</ID>21 </output>
<output>
<ID>OUT_3</ID>22 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>33</ID>
<type>DA_FROM</type>
<position>-28,-70.5</position>
<input>
<ID>IN_0</ID>269 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID MANUAL_DATA</lparam></gate>
<gate>
<ID>36</ID>
<type>DE_TO</type>
<position>93,-77.5</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A0</lparam></gate>
<gate>
<ID>37</ID>
<type>DE_TO</type>
<position>91,-77.5</position>
<input>
<ID>IN_0</ID>30 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A2</lparam></gate>
<gate>
<ID>38</ID>
<type>DE_TO</type>
<position>89,-77.5</position>
<input>
<ID>IN_0</ID>29 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A4</lparam></gate>
<gate>
<ID>39</ID>
<type>DE_TO</type>
<position>87,-77.5</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A6</lparam></gate>
<gate>
<ID>40</ID>
<type>DE_TO</type>
<position>92,-67</position>
<input>
<ID>IN_0</ID>35 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A1</lparam></gate>
<gate>
<ID>41</ID>
<type>DE_TO</type>
<position>90,-67</position>
<input>
<ID>IN_0</ID>36 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A3</lparam></gate>
<gate>
<ID>42</ID>
<type>DE_TO</type>
<position>88,-67</position>
<input>
<ID>IN_0</ID>37 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A5</lparam></gate>
<gate>
<ID>43</ID>
<type>BE_COMPARATOR_4BIT</type>
<position>77,-100.5</position>
<output>
<ID>A_equal_B</ID>49 </output>
<output>
<ID>A_greater_B</ID>47 </output>
<output>
<ID>A_less_B</ID>48 </output>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_2</ID>73 </input>
<input>
<ID>IN_3</ID>74 </input>
<input>
<ID>IN_B_0</ID>55 </input>
<input>
<ID>IN_B_1</ID>56 </input>
<input>
<ID>IN_B_2</ID>57 </input>
<input>
<ID>IN_B_3</ID>58 </input>
<input>
<ID>in_A_equal_B</ID>33 </input>
<input>
<ID>in_A_greater_B</ID>32 </input>
<input>
<ID>in_A_less_B</ID>34 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>44</ID>
<type>DE_TO</type>
<position>86,-67</position>
<input>
<ID>IN_0</ID>38 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A7</lparam></gate>
<gate>
<ID>45</ID>
<type>DE_TO</type>
<position>105,-77.5</position>
<input>
<ID>IN_0</ID>42 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B0</lparam></gate>
<gate>
<ID>46</ID>
<type>DE_TO</type>
<position>103,-77.5</position>
<input>
<ID>IN_0</ID>41 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B2</lparam></gate>
<gate>
<ID>47</ID>
<type>HA_JUNC_2</type>
<position>98,-80.5</position>
<input>
<ID>N_in0</ID>46 </input>
<input>
<ID>N_in1</ID>58 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>48</ID>
<type>HA_JUNC_2</type>
<position>99,-80.5</position>
<input>
<ID>N_in0</ID>39 </input>
<input>
<ID>N_in1</ID>57 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>49</ID>
<type>HA_JUNC_2</type>
<position>100,-80.5</position>
<input>
<ID>N_in0</ID>45 </input>
<input>
<ID>N_in1</ID>56 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>50</ID>
<type>HA_JUNC_2</type>
<position>101,-80.5</position>
<input>
<ID>N_in0</ID>40 </input>
<input>
<ID>N_in1</ID>55 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>51</ID>
<type>HA_JUNC_2</type>
<position>102,-80.5</position>
<input>
<ID>N_in0</ID>44 </input>
<input>
<ID>N_in1</ID>54 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>52</ID>
<type>AE_REGISTER8</type>
<position>30,5</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>65 </input>
<input>
<ID>IN_2</ID>59 </input>
<input>
<ID>IN_3</ID>63 </input>
<input>
<ID>IN_4</ID>62 </input>
<input>
<ID>IN_5</ID>60 </input>
<input>
<ID>IN_6</ID>64 </input>
<input>
<ID>IN_7</ID>66 </input>
<output>
<ID>OUT_0</ID>80 </output>
<output>
<ID>OUT_1</ID>81 </output>
<output>
<ID>OUT_2</ID>82 </output>
<output>
<ID>OUT_3</ID>83 </output>
<output>
<ID>OUT_4</ID>84 </output>
<output>
<ID>OUT_5</ID>85 </output>
<output>
<ID>OUT_6</ID>86 </output>
<output>
<ID>OUT_7</ID>87 </output>
<input>
<ID>clear</ID>77 </input>
<input>
<ID>clock</ID>156 </input>
<input>
<ID>load</ID>76 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 96</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>53</ID>
<type>HA_JUNC_2</type>
<position>103,-80.5</position>
<input>
<ID>N_in0</ID>41 </input>
<input>
<ID>N_in1</ID>53 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>54</ID>
<type>HA_JUNC_2</type>
<position>7,90.5</position>
<input>
<ID>N_in0</ID>120 </input>
<input>
<ID>N_in1</ID>66 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>55</ID>
<type>HA_JUNC_2</type>
<position>8,90.5</position>
<input>
<ID>N_in0</ID>116 </input>
<input>
<ID>N_in1</ID>64 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>56</ID>
<type>HA_JUNC_2</type>
<position>9,90.5</position>
<input>
<ID>N_in0</ID>119 </input>
<input>
<ID>N_in1</ID>60 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>57</ID>
<type>HA_JUNC_2</type>
<position>10,90.5</position>
<input>
<ID>N_in0</ID>115 </input>
<input>
<ID>N_in1</ID>62 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>58</ID>
<type>HA_JUNC_2</type>
<position>11,90.5</position>
<input>
<ID>N_in0</ID>118 </input>
<input>
<ID>N_in1</ID>63 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>59</ID>
<type>HA_JUNC_2</type>
<position>12,90.5</position>
<input>
<ID>N_in0</ID>113 </input>
<input>
<ID>N_in1</ID>59 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>60</ID>
<type>HA_JUNC_2</type>
<position>13,90.5</position>
<input>
<ID>N_in0</ID>117 </input>
<input>
<ID>N_in1</ID>65 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>61</ID>
<type>HA_JUNC_2</type>
<position>14,90.5</position>
<input>
<ID>N_in0</ID>114 </input>
<input>
<ID>N_in1</ID>61 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>62</ID>
<type>HA_JUNC_2</type>
<position>7,-121</position>
<input>
<ID>N_in0</ID>66 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>63</ID>
<type>HA_JUNC_2</type>
<position>8,-121</position>
<input>
<ID>N_in0</ID>64 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>64</ID>
<type>HA_JUNC_2</type>
<position>9,-121</position>
<input>
<ID>N_in0</ID>60 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>65</ID>
<type>HA_JUNC_2</type>
<position>10,-121</position>
<input>
<ID>N_in0</ID>62 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>66</ID>
<type>HA_JUNC_2</type>
<position>11,-121</position>
<input>
<ID>N_in0</ID>63 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>67</ID>
<type>HA_JUNC_2</type>
<position>12,-121</position>
<input>
<ID>N_in0</ID>59 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>68</ID>
<type>HA_JUNC_2</type>
<position>13,-121</position>
<input>
<ID>N_in0</ID>65 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>69</ID>
<type>HA_JUNC_2</type>
<position>14,-121</position>
<input>
<ID>N_in0</ID>61 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>70</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>86.5,12</position>
<input>
<ID>ENABLE_0</ID>79 </input>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>81 </input>
<input>
<ID>IN_2</ID>82 </input>
<input>
<ID>IN_3</ID>83 </input>
<input>
<ID>IN_4</ID>84 </input>
<input>
<ID>IN_5</ID>85 </input>
<input>
<ID>IN_6</ID>86 </input>
<input>
<ID>IN_7</ID>87 </input>
<output>
<ID>OUT_0</ID>99 </output>
<output>
<ID>OUT_1</ID>103 </output>
<output>
<ID>OUT_2</ID>100 </output>
<output>
<ID>OUT_3</ID>104 </output>
<output>
<ID>OUT_4</ID>101 </output>
<output>
<ID>OUT_5</ID>108 </output>
<output>
<ID>OUT_6</ID>102 </output>
<output>
<ID>OUT_7</ID>107 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>71</ID>
<type>HA_JUNC_2</type>
<position>104,-80.5</position>
<input>
<ID>N_in0</ID>43 </input>
<input>
<ID>N_in1</ID>52 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>72</ID>
<type>HA_JUNC_2</type>
<position>105,-80.5</position>
<input>
<ID>N_in0</ID>42 </input>
<input>
<ID>N_in1</ID>51 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>73</ID>
<type>HA_JUNC_2</type>
<position>86,-80.5</position>
<input>
<ID>N_in0</ID>38 </input>
<input>
<ID>N_in1</ID>74 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>30.5,17.5</position>
<gparam>LABEL_TEXT R16</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>HA_JUNC_2</type>
<position>87,-80.5</position>
<input>
<ID>N_in0</ID>28 </input>
<input>
<ID>N_in1</ID>73 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>76</ID>
<type>DA_FROM</type>
<position>26.5,12.5</position>
<input>
<ID>IN_0</ID>76 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R16_LD</lparam></gate>
<gate>
<ID>77</ID>
<type>DA_FROM</type>
<position>29,-3.5</position>
<input>
<ID>IN_0</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R16_CLR</lparam></gate>
<gate>
<ID>78</ID>
<type>DA_FROM</type>
<position>79.5,12</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R16_ALU_A</lparam></gate>
<gate>
<ID>79</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>110.5,12</position>
<input>
<ID>ENABLE_0</ID>88 </input>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>81 </input>
<input>
<ID>IN_2</ID>82 </input>
<input>
<ID>IN_3</ID>83 </input>
<input>
<ID>IN_4</ID>84 </input>
<input>
<ID>IN_5</ID>85 </input>
<input>
<ID>IN_6</ID>86 </input>
<input>
<ID>IN_7</ID>87 </input>
<output>
<ID>OUT_0</ID>110 </output>
<output>
<ID>OUT_1</ID>289 </output>
<output>
<ID>OUT_2</ID>109 </output>
<output>
<ID>OUT_3</ID>288 </output>
<output>
<ID>OUT_4</ID>111 </output>
<output>
<ID>OUT_5</ID>287 </output>
<output>
<ID>OUT_6</ID>112 </output>
<output>
<ID>OUT_7</ID>286 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>80</ID>
<type>DA_FROM</type>
<position>103.5,12</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R16_ALU_B</lparam></gate>
<gate>
<ID>81</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>62,12</position>
<input>
<ID>ENABLE_0</ID>89 </input>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>81 </input>
<input>
<ID>IN_2</ID>82 </input>
<input>
<ID>IN_3</ID>83 </input>
<input>
<ID>IN_4</ID>84 </input>
<input>
<ID>IN_5</ID>85 </input>
<input>
<ID>IN_6</ID>86 </input>
<input>
<ID>IN_7</ID>87 </input>
<output>
<ID>OUT_0</ID>90 </output>
<output>
<ID>OUT_1</ID>91 </output>
<output>
<ID>OUT_2</ID>92 </output>
<output>
<ID>OUT_3</ID>98 </output>
<output>
<ID>OUT_4</ID>93 </output>
<output>
<ID>OUT_5</ID>97 </output>
<output>
<ID>OUT_6</ID>94 </output>
<output>
<ID>OUT_7</ID>96 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>82</ID>
<type>DA_FROM</type>
<position>55,12</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R16_DATA</lparam></gate>
<gate>
<ID>83</ID>
<type>HA_JUNC_2</type>
<position>88,-80.5</position>
<input>
<ID>N_in0</ID>37 </input>
<input>
<ID>N_in1</ID>72 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>84</ID>
<type>HA_JUNC_2</type>
<position>89,-80.5</position>
<input>
<ID>N_in0</ID>29 </input>
<input>
<ID>N_in1</ID>71 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>85</ID>
<type>DE_TO</type>
<position>65.5,16</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>86</ID>
<type>DE_TO</type>
<position>64.5,21</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>87</ID>
<type>DE_TO</type>
<position>63.5,16</position>
<input>
<ID>IN_0</ID>92 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>88</ID>
<type>DE_TO</type>
<position>61.5,16</position>
<input>
<ID>IN_0</ID>93 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>89</ID>
<type>DE_TO</type>
<position>59.5,16</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>90</ID>
<type>HA_JUNC_2</type>
<position>90,-80.5</position>
<input>
<ID>N_in0</ID>36 </input>
<input>
<ID>N_in1</ID>70 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>91</ID>
<type>DE_TO</type>
<position>62.5,21</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>92</ID>
<type>DE_TO</type>
<position>60.5,21</position>
<input>
<ID>IN_0</ID>97 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>93</ID>
<type>DE_TO</type>
<position>58.5,21</position>
<input>
<ID>IN_0</ID>96 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>94</ID>
<type>DE_TO</type>
<position>90,16</position>
<input>
<ID>IN_0</ID>99 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A0</lparam></gate>
<gate>
<ID>95</ID>
<type>DE_TO</type>
<position>88,16</position>
<input>
<ID>IN_0</ID>100 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A2</lparam></gate>
<gate>
<ID>96</ID>
<type>DE_TO</type>
<position>86,16</position>
<input>
<ID>IN_0</ID>101 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A4</lparam></gate>
<gate>
<ID>97</ID>
<type>DE_TO</type>
<position>84,16</position>
<input>
<ID>IN_0</ID>102 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A6</lparam></gate>
<gate>
<ID>98</ID>
<type>DE_TO</type>
<position>89,26.5</position>
<input>
<ID>IN_0</ID>103 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A1</lparam></gate>
<gate>
<ID>99</ID>
<type>DE_TO</type>
<position>87,26.5</position>
<input>
<ID>IN_0</ID>104 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A3</lparam></gate>
<gate>
<ID>100</ID>
<type>DE_TO</type>
<position>85,26.5</position>
<input>
<ID>IN_0</ID>108 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A5</lparam></gate>
<gate>
<ID>101</ID>
<type>DE_TO</type>
<position>83,26.5</position>
<input>
<ID>IN_0</ID>107 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A7</lparam></gate>
<gate>
<ID>102</ID>
<type>DE_TO</type>
<position>114,16</position>
<input>
<ID>IN_0</ID>110 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B0</lparam></gate>
<gate>
<ID>103</ID>
<type>DE_TO</type>
<position>112,16</position>
<input>
<ID>IN_0</ID>109 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B2</lparam></gate>
<gate>
<ID>104</ID>
<type>DE_TO</type>
<position>110,16</position>
<input>
<ID>IN_0</ID>111 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B4</lparam></gate>
<gate>
<ID>105</ID>
<type>DE_TO</type>
<position>108,16</position>
<input>
<ID>IN_0</ID>112 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B6</lparam></gate>
<gate>
<ID>106</ID>
<type>DE_TO</type>
<position>113,26.5</position>
<input>
<ID>IN_0</ID>289 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B1</lparam></gate>
<gate>
<ID>107</ID>
<type>DE_TO</type>
<position>111,26.5</position>
<input>
<ID>IN_0</ID>288 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B3</lparam></gate>
<gate>
<ID>108</ID>
<type>DE_TO</type>
<position>109,26.5</position>
<input>
<ID>IN_0</ID>287 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B5</lparam></gate>
<gate>
<ID>109</ID>
<type>DE_TO</type>
<position>107,26.5</position>
<input>
<ID>IN_0</ID>286 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B7</lparam></gate>
<gate>
<ID>110</ID>
<type>DE_TO</type>
<position>14,93.5</position>
<input>
<ID>IN_0</ID>114 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>111</ID>
<type>DE_TO</type>
<position>13,98.5</position>
<input>
<ID>IN_0</ID>117 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>112</ID>
<type>DE_TO</type>
<position>12,93.5</position>
<input>
<ID>IN_0</ID>113 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>113</ID>
<type>DE_TO</type>
<position>10,93.5</position>
<input>
<ID>IN_0</ID>115 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>114</ID>
<type>DE_TO</type>
<position>8,93.5</position>
<input>
<ID>IN_0</ID>116 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>115</ID>
<type>DE_TO</type>
<position>11,98.5</position>
<input>
<ID>IN_0</ID>118 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>116</ID>
<type>DE_TO</type>
<position>9,98.5</position>
<input>
<ID>IN_0</ID>119 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>117</ID>
<type>DE_TO</type>
<position>7,98.5</position>
<input>
<ID>IN_0</ID>120 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>118</ID>
<type>HA_JUNC_2</type>
<position>91,-80.5</position>
<input>
<ID>N_in0</ID>30 </input>
<input>
<ID>N_in1</ID>69 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>119</ID>
<type>HA_JUNC_2</type>
<position>92,-80.5</position>
<input>
<ID>N_in0</ID>35 </input>
<input>
<ID>N_in1</ID>68 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>120</ID>
<type>HA_JUNC_2</type>
<position>93,-80.5</position>
<input>
<ID>N_in0</ID>31 </input>
<input>
<ID>N_in1</ID>67 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>121</ID>
<type>AE_REGISTER8</type>
<position>30,-33.5</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>65 </input>
<input>
<ID>IN_2</ID>59 </input>
<input>
<ID>IN_3</ID>63 </input>
<input>
<ID>IN_4</ID>62 </input>
<input>
<ID>IN_5</ID>60 </input>
<input>
<ID>IN_6</ID>64 </input>
<input>
<ID>IN_7</ID>66 </input>
<output>
<ID>OUT_0</ID>125 </output>
<output>
<ID>OUT_1</ID>126 </output>
<output>
<ID>OUT_2</ID>127 </output>
<output>
<ID>OUT_3</ID>128 </output>
<output>
<ID>OUT_4</ID>129 </output>
<output>
<ID>OUT_5</ID>130 </output>
<output>
<ID>OUT_6</ID>131 </output>
<output>
<ID>OUT_7</ID>132 </output>
<input>
<ID>clear</ID>123 </input>
<input>
<ID>clock</ID>155 </input>
<input>
<ID>load</ID>122 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>122</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>86.5,-26.5</position>
<input>
<ID>ENABLE_0</ID>124 </input>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>126 </input>
<input>
<ID>IN_2</ID>127 </input>
<input>
<ID>IN_3</ID>128 </input>
<input>
<ID>IN_4</ID>129 </input>
<input>
<ID>IN_5</ID>130 </input>
<input>
<ID>IN_6</ID>131 </input>
<input>
<ID>IN_7</ID>132 </input>
<output>
<ID>OUT_0</ID>143 </output>
<output>
<ID>OUT_1</ID>147 </output>
<output>
<ID>OUT_2</ID>144 </output>
<output>
<ID>OUT_3</ID>148 </output>
<output>
<ID>OUT_4</ID>145 </output>
<output>
<ID>OUT_5</ID>150 </output>
<output>
<ID>OUT_6</ID>146 </output>
<output>
<ID>OUT_7</ID>149 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_LABEL</type>
<position>30.5,-21</position>
<gparam>LABEL_TEXT R17</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>124</ID>
<type>DA_FROM</type>
<position>26.5,-26</position>
<input>
<ID>IN_0</ID>122 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R17_LD</lparam></gate>
<gate>
<ID>125</ID>
<type>DA_FROM</type>
<position>29,-41.5</position>
<input>
<ID>IN_0</ID>123 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R17_CLR</lparam></gate>
<gate>
<ID>126</ID>
<type>DA_FROM</type>
<position>79.5,-26.5</position>
<input>
<ID>IN_0</ID>124 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R17_ALU_A</lparam></gate>
<gate>
<ID>127</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>110.5,-26.5</position>
<input>
<ID>ENABLE_0</ID>133 </input>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>126 </input>
<input>
<ID>IN_2</ID>127 </input>
<input>
<ID>IN_3</ID>128 </input>
<input>
<ID>IN_4</ID>129 </input>
<input>
<ID>IN_5</ID>130 </input>
<input>
<ID>IN_6</ID>131 </input>
<input>
<ID>IN_7</ID>132 </input>
<output>
<ID>OUT_0</ID>152 </output>
<output>
<ID>OUT_1</ID>285 </output>
<output>
<ID>OUT_2</ID>151 </output>
<output>
<ID>OUT_3</ID>284 </output>
<output>
<ID>OUT_4</ID>153 </output>
<output>
<ID>OUT_5</ID>283 </output>
<output>
<ID>OUT_6</ID>154 </output>
<output>
<ID>OUT_7</ID>282 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>128</ID>
<type>DA_FROM</type>
<position>103.5,-26.5</position>
<input>
<ID>IN_0</ID>133 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R17_ALU_B</lparam></gate>
<gate>
<ID>129</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>62,-26.5</position>
<input>
<ID>ENABLE_0</ID>134 </input>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>126 </input>
<input>
<ID>IN_2</ID>127 </input>
<input>
<ID>IN_3</ID>128 </input>
<input>
<ID>IN_4</ID>129 </input>
<input>
<ID>IN_5</ID>130 </input>
<input>
<ID>IN_6</ID>131 </input>
<input>
<ID>IN_7</ID>132 </input>
<output>
<ID>OUT_0</ID>135 </output>
<output>
<ID>OUT_1</ID>136 </output>
<output>
<ID>OUT_2</ID>137 </output>
<output>
<ID>OUT_3</ID>142 </output>
<output>
<ID>OUT_4</ID>138 </output>
<output>
<ID>OUT_5</ID>141 </output>
<output>
<ID>OUT_6</ID>139 </output>
<output>
<ID>OUT_7</ID>140 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>130</ID>
<type>DA_FROM</type>
<position>55,-26.5</position>
<input>
<ID>IN_0</ID>134 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R17_DATA</lparam></gate>
<gate>
<ID>131</ID>
<type>DE_TO</type>
<position>65.5,-22.5</position>
<input>
<ID>IN_0</ID>135 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>132</ID>
<type>DE_TO</type>
<position>64.5,-17.5</position>
<input>
<ID>IN_0</ID>136 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>133</ID>
<type>DE_TO</type>
<position>63.5,-22.5</position>
<input>
<ID>IN_0</ID>137 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>134</ID>
<type>DE_TO</type>
<position>61.5,-22.5</position>
<input>
<ID>IN_0</ID>138 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>135</ID>
<type>DE_TO</type>
<position>59.5,-22.5</position>
<input>
<ID>IN_0</ID>139 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>136</ID>
<type>DE_TO</type>
<position>62.5,-17.5</position>
<input>
<ID>IN_0</ID>142 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>137</ID>
<type>DE_TO</type>
<position>60.5,-17.5</position>
<input>
<ID>IN_0</ID>141 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>138</ID>
<type>DE_TO</type>
<position>58.5,-17.5</position>
<input>
<ID>IN_0</ID>140 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>139</ID>
<type>DE_TO</type>
<position>90,-22.5</position>
<input>
<ID>IN_0</ID>143 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A0</lparam></gate>
<gate>
<ID>140</ID>
<type>DE_TO</type>
<position>88,-22.5</position>
<input>
<ID>IN_0</ID>144 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A2</lparam></gate>
<gate>
<ID>141</ID>
<type>DE_TO</type>
<position>86,-22.5</position>
<input>
<ID>IN_0</ID>145 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A4</lparam></gate>
<gate>
<ID>142</ID>
<type>DE_TO</type>
<position>84,-22.5</position>
<input>
<ID>IN_0</ID>146 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A6</lparam></gate>
<gate>
<ID>143</ID>
<type>DE_TO</type>
<position>89,-12</position>
<input>
<ID>IN_0</ID>147 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A1</lparam></gate>
<gate>
<ID>144</ID>
<type>DE_TO</type>
<position>87,-12</position>
<input>
<ID>IN_0</ID>148 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A3</lparam></gate>
<gate>
<ID>145</ID>
<type>DE_TO</type>
<position>85,-12</position>
<input>
<ID>IN_0</ID>150 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A5</lparam></gate>
<gate>
<ID>146</ID>
<type>DE_TO</type>
<position>83,-12</position>
<input>
<ID>IN_0</ID>149 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A7</lparam></gate>
<gate>
<ID>147</ID>
<type>DE_TO</type>
<position>114,-22.5</position>
<input>
<ID>IN_0</ID>152 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B0</lparam></gate>
<gate>
<ID>148</ID>
<type>DE_TO</type>
<position>112,-22.5</position>
<input>
<ID>IN_0</ID>151 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B2</lparam></gate>
<gate>
<ID>149</ID>
<type>DE_TO</type>
<position>110,-22.5</position>
<input>
<ID>IN_0</ID>153 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B4</lparam></gate>
<gate>
<ID>150</ID>
<type>DE_TO</type>
<position>108,-22.5</position>
<input>
<ID>IN_0</ID>154 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B6</lparam></gate>
<gate>
<ID>151</ID>
<type>DE_TO</type>
<position>113,-12</position>
<input>
<ID>IN_0</ID>285 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B1</lparam></gate>
<gate>
<ID>152</ID>
<type>DE_TO</type>
<position>111,-12</position>
<input>
<ID>IN_0</ID>284 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B3</lparam></gate>
<gate>
<ID>153</ID>
<type>DE_TO</type>
<position>109,-12</position>
<input>
<ID>IN_0</ID>283 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B5</lparam></gate>
<gate>
<ID>154</ID>
<type>DE_TO</type>
<position>107,-12</position>
<input>
<ID>IN_0</ID>282 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B7</lparam></gate>
<gate>
<ID>155</ID>
<type>DA_FROM</type>
<position>27,-39.5</position>
<input>
<ID>IN_0</ID>155 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>156</ID>
<type>DA_FROM</type>
<position>27,-1</position>
<input>
<ID>IN_0</ID>156 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>157</ID>
<type>DA_FROM</type>
<position>-26,-7.5</position>
<input>
<ID>IN_0</ID>157 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID CLK</lparam></gate>
<gate>
<ID>158</ID>
<type>DE_TO</type>
<position>101,-77.5</position>
<input>
<ID>IN_0</ID>40 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B4</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_TOGGLE</type>
<position>-30,-7.5</position>
<output>
<ID>OUT_0</ID>157 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>160</ID>
<type>DE_TO</type>
<position>99,-77.5</position>
<input>
<ID>IN_0</ID>39 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B6</lparam></gate>
<gate>
<ID>161</ID>
<type>DE_TO</type>
<position>104,-67</position>
<input>
<ID>IN_0</ID>43 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B1</lparam></gate>
<gate>
<ID>162</ID>
<type>DE_TO</type>
<position>102,-67</position>
<input>
<ID>IN_0</ID>44 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B3</lparam></gate>
<gate>
<ID>163</ID>
<type>DE_TO</type>
<position>100,-67</position>
<input>
<ID>IN_0</ID>45 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B5</lparam></gate>
<gate>
<ID>164</ID>
<type>DE_TO</type>
<position>98,-67</position>
<input>
<ID>IN_0</ID>46 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B7</lparam></gate>
<gate>
<ID>165</ID>
<type>DE_TO</type>
<position>67,-98.5</position>
<input>
<ID>IN_0</ID>47 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID ALU_A_GREATER</lparam></gate>
<gate>
<ID>166</ID>
<type>DE_TO</type>
<position>67,-102.5</position>
<input>
<ID>IN_0</ID>48 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID ALU_A_LESS</lparam></gate>
<gate>
<ID>167</ID>
<type>DE_TO</type>
<position>67,-100.5</position>
<input>
<ID>IN_0</ID>49 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID ALU_EQUAL</lparam></gate>
<gate>
<ID>168</ID>
<type>DE_TO</type>
<position>98.5,-105.5</position>
<input>
<ID>IN_0</ID>50 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID ALU_CARRY_OUT</lparam></gate>
<gate>
<ID>169</ID>
<type>DE_TO</type>
<position>138,-99</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ALU_CARRY_IN</lparam></gate>
<gate>
<ID>170</ID>
<type>DE_TO</type>
<position>98.5,-108</position>
<input>
<ID>IN_0</ID>78 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID ALU_SIGNED_CARRY_OUT</lparam></gate>
<gate>
<ID>171</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>120,-116</position>
<input>
<ID>ENABLE_0</ID>95 </input>
<input>
<ID>IN_0</ID>163 </input>
<input>
<ID>IN_1</ID>164 </input>
<input>
<ID>IN_2</ID>165 </input>
<input>
<ID>IN_3</ID>166 </input>
<input>
<ID>IN_4</ID>167 </input>
<input>
<ID>IN_5</ID>168 </input>
<input>
<ID>IN_6</ID>169 </input>
<input>
<ID>IN_7</ID>170 </input>
<output>
<ID>OUT_0</ID>105 </output>
<output>
<ID>OUT_1</ID>106 </output>
<output>
<ID>OUT_2</ID>121 </output>
<output>
<ID>OUT_3</ID>162 </output>
<output>
<ID>OUT_4</ID>158 </output>
<output>
<ID>OUT_5</ID>161 </output>
<output>
<ID>OUT_6</ID>159 </output>
<output>
<ID>OUT_7</ID>160 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>172</ID>
<type>DA_FROM</type>
<position>109,-116</position>
<input>
<ID>IN_0</ID>95 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ALU_DATA</lparam></gate>
<gate>
<ID>173</ID>
<type>DE_TO</type>
<position>123.5,-112</position>
<input>
<ID>IN_0</ID>105 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>174</ID>
<type>DE_TO</type>
<position>122.5,-107</position>
<input>
<ID>IN_0</ID>106 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>175</ID>
<type>DE_TO</type>
<position>121.5,-112</position>
<input>
<ID>IN_0</ID>121 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>176</ID>
<type>DE_TO</type>
<position>119.5,-112</position>
<input>
<ID>IN_0</ID>158 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>177</ID>
<type>DE_TO</type>
<position>117.5,-112</position>
<input>
<ID>IN_0</ID>159 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>178</ID>
<type>DE_TO</type>
<position>120.5,-107</position>
<input>
<ID>IN_0</ID>162 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>179</ID>
<type>DE_TO</type>
<position>118.5,-107</position>
<input>
<ID>IN_0</ID>161 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>180</ID>
<type>DE_TO</type>
<position>116.5,-107</position>
<input>
<ID>IN_0</ID>160 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>190</ID>
<type>DE_TO</type>
<position>32.5,-69.5</position>
<input>
<ID>IN_0</ID>182 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A0</lparam></gate>
<gate>
<ID>191</ID>
<type>DE_TO</type>
<position>30.5,-69.5</position>
<input>
<ID>IN_0</ID>181 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A2</lparam></gate>
<gate>
<ID>192</ID>
<type>DE_TO</type>
<position>28.5,-69.5</position>
<input>
<ID>IN_0</ID>180 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A4</lparam></gate>
<gate>
<ID>193</ID>
<type>DE_TO</type>
<position>26.5,-69.5</position>
<input>
<ID>IN_0</ID>179 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A6</lparam></gate>
<gate>
<ID>194</ID>
<type>DE_TO</type>
<position>31.5,-59</position>
<input>
<ID>IN_0</ID>183 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A1</lparam></gate>
<gate>
<ID>195</ID>
<type>DE_TO</type>
<position>29.5,-59</position>
<input>
<ID>IN_0</ID>184 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A3</lparam></gate>
<gate>
<ID>196</ID>
<type>DE_TO</type>
<position>27.5,-59</position>
<input>
<ID>IN_0</ID>185 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A5</lparam></gate>
<gate>
<ID>197</ID>
<type>DE_TO</type>
<position>25.5,-59</position>
<input>
<ID>IN_0</ID>186 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_A7</lparam></gate>
<gate>
<ID>198</ID>
<type>DE_TO</type>
<position>50.5,-69.5</position>
<input>
<ID>IN_0</ID>190 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B0</lparam></gate>
<gate>
<ID>199</ID>
<type>DE_TO</type>
<position>48.5,-69.5</position>
<input>
<ID>IN_0</ID>189 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B2</lparam></gate>
<gate>
<ID>200</ID>
<type>HA_JUNC_2</type>
<position>43.5,-72.5</position>
<input>
<ID>N_in0</ID>194 </input>
<input>
<ID>N_in1</ID>196 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>201</ID>
<type>HA_JUNC_2</type>
<position>44.5,-72.5</position>
<input>
<ID>N_in0</ID>187 </input>
<input>
<ID>N_in1</ID>197 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>202</ID>
<type>HA_JUNC_2</type>
<position>45.5,-72.5</position>
<input>
<ID>N_in0</ID>193 </input>
<input>
<ID>N_in1</ID>200 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>203</ID>
<type>HA_JUNC_2</type>
<position>46.5,-72.5</position>
<input>
<ID>N_in0</ID>188 </input>
<input>
<ID>N_in1</ID>201 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>204</ID>
<type>HA_JUNC_2</type>
<position>47.5,-72.5</position>
<input>
<ID>N_in0</ID>192 </input>
<input>
<ID>N_in1</ID>198 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>205</ID>
<type>HA_JUNC_2</type>
<position>48.5,-72.5</position>
<input>
<ID>N_in0</ID>189 </input>
<input>
<ID>N_in1</ID>202 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>206</ID>
<type>HA_JUNC_2</type>
<position>49.5,-72.5</position>
<input>
<ID>N_in0</ID>191 </input>
<input>
<ID>N_in1</ID>199 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>207</ID>
<type>HA_JUNC_2</type>
<position>50.5,-72.5</position>
<input>
<ID>N_in0</ID>190 </input>
<input>
<ID>N_in1</ID>195 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>208</ID>
<type>HA_JUNC_2</type>
<position>25.5,-72.5</position>
<input>
<ID>N_in0</ID>186 </input>
<input>
<ID>N_in1</ID>203 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>209</ID>
<type>HA_JUNC_2</type>
<position>26.5,-72.5</position>
<input>
<ID>N_in0</ID>179 </input>
<input>
<ID>N_in1</ID>210 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>210</ID>
<type>HA_JUNC_2</type>
<position>27.5,-72.5</position>
<input>
<ID>N_in0</ID>185 </input>
<input>
<ID>N_in1</ID>204 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>211</ID>
<type>HA_JUNC_2</type>
<position>28.5,-72.5</position>
<input>
<ID>N_in0</ID>180 </input>
<input>
<ID>N_in1</ID>205 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>212</ID>
<type>HA_JUNC_2</type>
<position>29.5,-72.5</position>
<input>
<ID>N_in0</ID>184 </input>
<input>
<ID>N_in1</ID>206 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>213</ID>
<type>HA_JUNC_2</type>
<position>30.5,-72.5</position>
<input>
<ID>N_in0</ID>181 </input>
<input>
<ID>N_in1</ID>207 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>214</ID>
<type>HA_JUNC_2</type>
<position>31.5,-72.5</position>
<input>
<ID>N_in0</ID>183 </input>
<input>
<ID>N_in1</ID>209 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>215</ID>
<type>HA_JUNC_2</type>
<position>32.5,-72.5</position>
<input>
<ID>N_in0</ID>182 </input>
<input>
<ID>N_in1</ID>208 </input>
<gparam>LED_BOX -0.25,-0.25,0.25,0.25</gparam>
<gparam>angle 270</gparam></gate>
<gate>
<ID>216</ID>
<type>DE_TO</type>
<position>46.5,-69.5</position>
<input>
<ID>IN_0</ID>188 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B4</lparam></gate>
<gate>
<ID>217</ID>
<type>DE_TO</type>
<position>44.5,-69.5</position>
<input>
<ID>IN_0</ID>187 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B6</lparam></gate>
<gate>
<ID>218</ID>
<type>DE_TO</type>
<position>49.5,-59</position>
<input>
<ID>IN_0</ID>191 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B1</lparam></gate>
<gate>
<ID>219</ID>
<type>DE_TO</type>
<position>47.5,-59</position>
<input>
<ID>IN_0</ID>192 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B3</lparam></gate>
<gate>
<ID>220</ID>
<type>DE_TO</type>
<position>45.5,-59</position>
<input>
<ID>IN_0</ID>193 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B5</lparam></gate>
<gate>
<ID>221</ID>
<type>DE_TO</type>
<position>43.5,-59</position>
<input>
<ID>IN_0</ID>194 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_B7</lparam></gate>
<gate>
<ID>223</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>47,-75.5</position>
<input>
<ID>ENABLE_0</ID>211 </input>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>65 </input>
<input>
<ID>IN_2</ID>59 </input>
<input>
<ID>IN_3</ID>63 </input>
<input>
<ID>IN_4</ID>62 </input>
<input>
<ID>IN_5</ID>60 </input>
<input>
<ID>IN_6</ID>64 </input>
<input>
<ID>IN_7</ID>66 </input>
<output>
<ID>OUT_0</ID>195 </output>
<output>
<ID>OUT_1</ID>199 </output>
<output>
<ID>OUT_2</ID>202 </output>
<output>
<ID>OUT_3</ID>198 </output>
<output>
<ID>OUT_4</ID>201 </output>
<output>
<ID>OUT_5</ID>200 </output>
<output>
<ID>OUT_6</ID>197 </output>
<output>
<ID>OUT_7</ID>196 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>224</ID>
<type>BO_TRI_STATE_8BIT</type>
<position>29,-75.5</position>
<input>
<ID>ENABLE_0</ID>212 </input>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>65 </input>
<input>
<ID>IN_2</ID>59 </input>
<input>
<ID>IN_3</ID>63 </input>
<input>
<ID>IN_4</ID>62 </input>
<input>
<ID>IN_5</ID>60 </input>
<input>
<ID>IN_6</ID>64 </input>
<input>
<ID>IN_7</ID>66 </input>
<output>
<ID>OUT_0</ID>208 </output>
<output>
<ID>OUT_1</ID>209 </output>
<output>
<ID>OUT_2</ID>207 </output>
<output>
<ID>OUT_3</ID>206 </output>
<output>
<ID>OUT_4</ID>205 </output>
<output>
<ID>OUT_5</ID>204 </output>
<output>
<ID>OUT_6</ID>210 </output>
<output>
<ID>OUT_7</ID>203 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>225</ID>
<type>DE_TO</type>
<position>41,-72.5</position>
<input>
<ID>IN_0</ID>211 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_DATA_B</lparam></gate>
<gate>
<ID>226</ID>
<type>DE_TO</type>
<position>23,-72.5</position>
<input>
<ID>IN_0</ID>212 </input>
<gparam>angle 90</gparam>
<lparam>JUNCTION_ID ALU_DATA_A</lparam></gate>
<gate>
<ID>231</ID>
<type>DA_FROM</type>
<position>-28,-87.5</position>
<input>
<ID>IN_0</ID>237 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID ALU_DATA</lparam></gate>
<gate>
<ID>234</ID>
<type>BI_DECODER_4x16</type>
<position>-33,-63</position>
<input>
<ID>ENABLE</ID>230 </input>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>219 </input>
<input>
<ID>IN_2</ID>220 </input>
<input>
<ID>IN_3</ID>221 </input>
<output>
<ID>OUT_0</ID>269 </output>
<output>
<ID>OUT_15</ID>239 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>235</ID>
<type>BI_DECODER_4x16</type>
<position>-33,-80</position>
<input>
<ID>ENABLE</ID>229 </input>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>219 </input>
<input>
<ID>IN_2</ID>220 </input>
<input>
<ID>IN_3</ID>221 </input>
<output>
<ID>OUT_0</ID>237 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>241</ID>
<type>DD_KEYPAD_HEX</type>
<position>-57,-70.5</position>
<output>
<ID>OUT_0</ID>218 </output>
<output>
<ID>OUT_1</ID>219 </output>
<output>
<ID>OUT_2</ID>220 </output>
<output>
<ID>OUT_3</ID>221 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>242</ID>
<type>DD_KEYPAD_HEX</type>
<position>-69,-70.5</position>
<output>
<ID>OUT_0</ID>224 </output>
<output>
<ID>OUT_1</ID>225 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>244</ID>
<type>BA_DECODER_2x4</type>
<position>-58.5,-84</position>
<input>
<ID>ENABLE</ID>226 </input>
<input>
<ID>IN_0</ID>224 </input>
<input>
<ID>IN_1</ID>225 </input>
<output>
<ID>OUT_0</ID>227 </output>
<output>
<ID>OUT_1</ID>228 </output>
<output>
<ID>OUT_2</ID>229 </output>
<output>
<ID>OUT_3</ID>230 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>246</ID>
<type>EE_VDD</type>
<position>-62,-81</position>
<output>
<ID>OUT_0</ID>226 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>247</ID>
<type>BI_DECODER_4x16</type>
<position>-33,-97</position>
<input>
<ID>ENABLE</ID>228 </input>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>219 </input>
<input>
<ID>IN_2</ID>220 </input>
<input>
<ID>IN_3</ID>221 </input>
<output>
<ID>OUT_0</ID>240 </output>
<output>
<ID>OUT_1</ID>236 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>248</ID>
<type>BI_DECODER_4x16</type>
<position>-33,-114</position>
<input>
<ID>ENABLE</ID>227 </input>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>219 </input>
<input>
<ID>IN_2</ID>220 </input>
<input>
<ID>IN_3</ID>221 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>249</ID>
<type>DA_FROM</type>
<position>-28,-55.5</position>
<input>
<ID>IN_0</ID>239 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID DATA_BUS_RELEASED</lparam></gate>
<gate>
<ID>251</ID>
<type>AA_LABEL</type>
<position>-82,-58</position>
<gparam>LABEL_TEXT DATA BUS SOURCE SELECTOR</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>252</ID>
<type>AA_LABEL</type>
<position>173.5,-51</position>
<gparam>LABEL_TEXT ALU A CHANNEL SOURCE SELECTOR</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>253</ID>
<type>AA_LABEL</type>
<position>261.5,-49.5</position>
<gparam>LABEL_TEXT ALU B CHANNEL SOURCE SELECTOR</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>254</ID>
<type>BI_DECODER_4x16</type>
<position>206,-62.5</position>
<input>
<ID>ENABLE</ID>251 </input>
<input>
<ID>IN_0</ID>241 </input>
<input>
<ID>IN_1</ID>242 </input>
<input>
<ID>IN_2</ID>243 </input>
<input>
<ID>IN_3</ID>244 </input>
<output>
<ID>OUT_0</ID>268 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>255</ID>
<type>BI_DECODER_4x16</type>
<position>206,-79.5</position>
<input>
<ID>ENABLE</ID>250 </input>
<input>
<ID>IN_0</ID>241 </input>
<input>
<ID>IN_1</ID>242 </input>
<input>
<ID>IN_2</ID>243 </input>
<input>
<ID>IN_3</ID>244 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>256</ID>
<type>DD_KEYPAD_HEX</type>
<position>182,-70</position>
<output>
<ID>OUT_0</ID>241 </output>
<output>
<ID>OUT_1</ID>242 </output>
<output>
<ID>OUT_2</ID>243 </output>
<output>
<ID>OUT_3</ID>244 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>257</ID>
<type>DD_KEYPAD_HEX</type>
<position>170,-70</position>
<output>
<ID>OUT_0</ID>245 </output>
<output>
<ID>OUT_1</ID>246 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>258</ID>
<type>BA_DECODER_2x4</type>
<position>180.5,-83.5</position>
<input>
<ID>ENABLE</ID>247 </input>
<input>
<ID>IN_0</ID>245 </input>
<input>
<ID>IN_1</ID>246 </input>
<output>
<ID>OUT_0</ID>248 </output>
<output>
<ID>OUT_1</ID>249 </output>
<output>
<ID>OUT_2</ID>250 </output>
<output>
<ID>OUT_3</ID>251 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>259</ID>
<type>EE_VDD</type>
<position>177,-80.5</position>
<output>
<ID>OUT_0</ID>247 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>260</ID>
<type>BI_DECODER_4x16</type>
<position>206,-96.5</position>
<input>
<ID>ENABLE</ID>249 </input>
<input>
<ID>IN_0</ID>241 </input>
<input>
<ID>IN_1</ID>242 </input>
<input>
<ID>IN_2</ID>243 </input>
<input>
<ID>IN_3</ID>244 </input>
<output>
<ID>OUT_0</ID>263 </output>
<output>
<ID>OUT_1</ID>264 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>261</ID>
<type>BI_DECODER_4x16</type>
<position>206,-113.5</position>
<input>
<ID>ENABLE</ID>248 </input>
<input>
<ID>IN_0</ID>241 </input>
<input>
<ID>IN_1</ID>242 </input>
<input>
<ID>IN_2</ID>243 </input>
<input>
<ID>IN_3</ID>244 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>262</ID>
<type>BI_DECODER_4x16</type>
<position>274.5,-61.5</position>
<input>
<ID>ENABLE</ID>262 </input>
<input>
<ID>IN_0</ID>252 </input>
<input>
<ID>IN_1</ID>253 </input>
<input>
<ID>IN_2</ID>254 </input>
<input>
<ID>IN_3</ID>255 </input>
<output>
<ID>OUT_0</ID>267 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>263</ID>
<type>BI_DECODER_4x16</type>
<position>274.5,-78.5</position>
<input>
<ID>ENABLE</ID>261 </input>
<input>
<ID>IN_0</ID>252 </input>
<input>
<ID>IN_1</ID>253 </input>
<input>
<ID>IN_2</ID>254 </input>
<input>
<ID>IN_3</ID>255 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>264</ID>
<type>DD_KEYPAD_HEX</type>
<position>250.5,-69</position>
<output>
<ID>OUT_0</ID>252 </output>
<output>
<ID>OUT_1</ID>253 </output>
<output>
<ID>OUT_2</ID>254 </output>
<output>
<ID>OUT_3</ID>255 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>265</ID>
<type>DD_KEYPAD_HEX</type>
<position>238.5,-69</position>
<output>
<ID>OUT_0</ID>256 </output>
<output>
<ID>OUT_1</ID>257 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>266</ID>
<type>BA_DECODER_2x4</type>
<position>249,-82.5</position>
<input>
<ID>ENABLE</ID>258 </input>
<input>
<ID>IN_0</ID>256 </input>
<input>
<ID>IN_1</ID>257 </input>
<output>
<ID>OUT_0</ID>259 </output>
<output>
<ID>OUT_1</ID>260 </output>
<output>
<ID>OUT_2</ID>261 </output>
<output>
<ID>OUT_3</ID>262 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>267</ID>
<type>EE_VDD</type>
<position>245.5,-79.5</position>
<output>
<ID>OUT_0</ID>258 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>268</ID>
<type>BI_DECODER_4x16</type>
<position>274.5,-95.5</position>
<input>
<ID>ENABLE</ID>260 </input>
<input>
<ID>IN_0</ID>252 </input>
<input>
<ID>IN_1</ID>253 </input>
<input>
<ID>IN_2</ID>254 </input>
<input>
<ID>IN_3</ID>255 </input>
<output>
<ID>OUT_0</ID>265 </output>
<output>
<ID>OUT_1</ID>266 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>269</ID>
<type>BI_DECODER_4x16</type>
<position>274.5,-112.5</position>
<input>
<ID>ENABLE</ID>259 </input>
<input>
<ID>IN_0</ID>252 </input>
<input>
<ID>IN_1</ID>253 </input>
<input>
<ID>IN_2</ID>254 </input>
<input>
<ID>IN_3</ID>255 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>270</ID>
<type>DA_FROM</type>
<position>211,-104</position>
<input>
<ID>IN_0</ID>263 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID R16_ALU_A</lparam></gate>
<gate>
<ID>271</ID>
<type>DA_FROM</type>
<position>226,-103</position>
<input>
<ID>IN_0</ID>264 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID R17_ALU_A</lparam></gate>
<gate>
<ID>272</ID>
<type>DA_FROM</type>
<position>279.5,-103</position>
<input>
<ID>IN_0</ID>265 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID R16_ALU_B</lparam></gate>
<gate>
<ID>273</ID>
<type>DA_FROM</type>
<position>294,-102</position>
<input>
<ID>IN_0</ID>266 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID R17_ALU_B</lparam></gate>
<gate>
<ID>274</ID>
<type>DE_TO</type>
<position>279.5,-69</position>
<input>
<ID>IN_0</ID>267 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ALU_DATA_B</lparam></gate>
<gate>
<ID>275</ID>
<type>DE_TO</type>
<position>211,-70</position>
<input>
<ID>IN_0</ID>268 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ALU_DATA_A</lparam></gate>
<gate>
<ID>277</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>-69.5,-23.5</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>278 </input>
<input>
<ID>IN_2</ID>272 </input>
<input>
<ID>IN_3</ID>277 </input>
<input>
<ID>IN_4</ID>273 </input>
<input>
<ID>IN_5</ID>276 </input>
<input>
<ID>IN_6</ID>274 </input>
<input>
<ID>IN_7</ID>275 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 98</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>278</ID>
<type>DE_TO</type>
<position>-76.5,-26.5</position>
<input>
<ID>IN_0</ID>270 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>279</ID>
<type>DE_TO</type>
<position>-82,-25.5</position>
<input>
<ID>IN_0</ID>278 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>280</ID>
<type>DE_TO</type>
<position>-76.5,-24.5</position>
<input>
<ID>IN_0</ID>272 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>281</ID>
<type>DE_TO</type>
<position>-76.5,-22.5</position>
<input>
<ID>IN_0</ID>273 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>282</ID>
<type>DE_TO</type>
<position>-76.5,-20.5</position>
<input>
<ID>IN_0</ID>274 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>283</ID>
<type>DE_TO</type>
<position>-82,-23.5</position>
<input>
<ID>IN_0</ID>277 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>284</ID>
<type>DE_TO</type>
<position>-82,-21.5</position>
<input>
<ID>IN_0</ID>276 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>285</ID>
<type>DE_TO</type>
<position>-82,-19.5</position>
<input>
<ID>IN_0</ID>275 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>286</ID>
<type>DE_TO</type>
<position>-26,-24.5</position>
<input>
<ID>IN_0</ID>279 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ALU_CARRY_IN</lparam></gate>
<gate>
<ID>287</ID>
<type>AA_TOGGLE</type>
<position>-30,-24.5</position>
<output>
<ID>OUT_0</ID>279 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>288</ID>
<type>DA_FROM</type>
<position>-26,-29</position>
<input>
<ID>IN_0</ID>280 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID R16_CLR</lparam></gate>
<gate>
<ID>289</ID>
<type>DA_FROM</type>
<position>-26,-32</position>
<input>
<ID>IN_0</ID>281 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID R17_CLR</lparam></gate>
<gate>
<ID>290</ID>
<type>AA_TOGGLE</type>
<position>-30,-29</position>
<output>
<ID>OUT_0</ID>280 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>291</ID>
<type>AA_TOGGLE</type>
<position>-30,-32</position>
<output>
<ID>OUT_0</ID>281 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>292</ID>
<type>DE_TO</type>
<position>123,-80</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 0</gparam>
<lparam>JUNCTION_ID ALU_HALF_CARRY_OUT</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-17,-28,-17</points>
<connection>
<GID>1</GID>
<name>IN_0</name></connection>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-20,-28,-20</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>3</ID>
<points>120,-99,120,-80</points>
<connection>
<GID>25</GID>
<name>carry_out</name></connection>
<connection>
<GID>24</GID>
<name>carry_in</name></connection>
<intersection>-80 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>120,-80,121,-80</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<intersection>120 3</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-36.5,15.5,-36.5,15.5</points>
<connection>
<GID>17</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>18</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,17.5,-28,17.5</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<connection>
<GID>19</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,17.5,-29,22.5</points>
<connection>
<GID>17</GID>
<name>OUT_1</name></connection>
<connection>
<GID>20</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,17.5,-30,17.5</points>
<connection>
<GID>17</GID>
<name>OUT_2</name></connection>
<connection>
<GID>21</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32,17.5,-32,17.5</points>
<connection>
<GID>17</GID>
<name>OUT_4</name></connection>
<connection>
<GID>23</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,17.5,-34,17.5</points>
<connection>
<GID>17</GID>
<name>OUT_6</name></connection>
<connection>
<GID>26</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,17.5,-35,22.5</points>
<connection>
<GID>17</GID>
<name>OUT_7</name></connection>
<connection>
<GID>29</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33,17.5,-33,22.5</points>
<connection>
<GID>17</GID>
<name>OUT_5</name></connection>
<connection>
<GID>28</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31,17.5,-31,22.5</points>
<connection>
<GID>17</GID>
<name>OUT_3</name></connection>
<connection>
<GID>27</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,5,-28,13.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48.5,5,-28,5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>-28 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,7,-29,13.5</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48.5,7,-29,7</points>
<connection>
<GID>32</GID>
<name>OUT_1</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,9,-30,13.5</points>
<connection>
<GID>17</GID>
<name>IN_2</name></connection>
<intersection>9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48.5,9,-30,9</points>
<connection>
<GID>32</GID>
<name>OUT_2</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31,11,-31,13.5</points>
<connection>
<GID>17</GID>
<name>IN_3</name></connection>
<intersection>11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-48.5,11,-31,11</points>
<connection>
<GID>32</GID>
<name>OUT_3</name></connection>
<intersection>-31 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32,0,-32,13.5</points>
<connection>
<GID>17</GID>
<name>IN_4</name></connection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-60,0,-32,0</points>
<intersection>-60 2</intersection>
<intersection>-32 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-60,0,-60,5</points>
<intersection>0 1</intersection>
<intersection>5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-60.5,5,-60,5</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>-60 2</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33,0.5,-33,13.5</points>
<connection>
<GID>17</GID>
<name>IN_5</name></connection>
<intersection>0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-59.5,0.5,-33,0.5</points>
<intersection>-59.5 2</intersection>
<intersection>-33 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-59.5,0.5,-59.5,7</points>
<intersection>0.5 1</intersection>
<intersection>7 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-60.5,7,-59.5,7</points>
<connection>
<GID>31</GID>
<name>OUT_1</name></connection>
<intersection>-59.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-34,1,-34,13.5</points>
<connection>
<GID>17</GID>
<name>IN_6</name></connection>
<intersection>1 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-59,1,-34,1</points>
<intersection>-59 2</intersection>
<intersection>-34 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-59,1,-59,9</points>
<intersection>1 1</intersection>
<intersection>9 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-60.5,9,-59,9</points>
<connection>
<GID>31</GID>
<name>OUT_2</name></connection>
<intersection>-59 2</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-35,1.5,-35,13.5</points>
<connection>
<GID>17</GID>
<name>IN_7</name></connection>
<intersection>1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-58.5,1.5,-35,1.5</points>
<intersection>-58.5 2</intersection>
<intersection>-35 0</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-58.5,1.5,-58.5,11</points>
<intersection>1.5 1</intersection>
<intersection>11 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-60.5,11,-58.5,11</points>
<connection>
<GID>31</GID>
<name>OUT_3</name></connection>
<intersection>-58.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-79.5,87,-79.5</points>
<connection>
<GID>75</GID>
<name>N_in0</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-79.5,89,-79.5</points>
<connection>
<GID>84</GID>
<name>N_in0</name></connection>
<connection>
<GID>38</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-79.5,91,-79.5</points>
<connection>
<GID>118</GID>
<name>N_in0</name></connection>
<connection>
<GID>37</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-79.5,93,-79.5</points>
<connection>
<GID>120</GID>
<name>N_in0</name></connection>
<connection>
<GID>36</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>85,-98.5,85,-98.5</points>
<connection>
<GID>22</GID>
<name>A_greater_B</name></connection>
<connection>
<GID>43</GID>
<name>in_A_greater_B</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>85,-100.5,85,-100.5</points>
<connection>
<GID>22</GID>
<name>A_equal_B</name></connection>
<connection>
<GID>43</GID>
<name>in_A_equal_B</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>85,-102.5,85,-102.5</points>
<connection>
<GID>22</GID>
<name>A_less_B</name></connection>
<connection>
<GID>43</GID>
<name>in_A_less_B</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,-79.5,92,-69</points>
<connection>
<GID>119</GID>
<name>N_in0</name></connection>
<connection>
<GID>40</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-79.5,90,-69</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<connection>
<GID>90</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-79.5,88,-69</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<connection>
<GID>83</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-79.5,86,-69</points>
<connection>
<GID>73</GID>
<name>N_in0</name></connection>
<connection>
<GID>44</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-79.5,99,-79.5</points>
<connection>
<GID>48</GID>
<name>N_in0</name></connection>
<connection>
<GID>160</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>101,-79.5,101,-79.5</points>
<connection>
<GID>50</GID>
<name>N_in0</name></connection>
<connection>
<GID>158</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-79.5,103,-79.5</points>
<connection>
<GID>53</GID>
<name>N_in0</name></connection>
<connection>
<GID>46</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-79.5,105,-79.5</points>
<connection>
<GID>72</GID>
<name>N_in0</name></connection>
<connection>
<GID>45</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-79.5,104,-69</points>
<connection>
<GID>71</GID>
<name>N_in0</name></connection>
<connection>
<GID>161</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-79.5,102,-69</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<connection>
<GID>51</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-79.5,100,-69</points>
<connection>
<GID>49</GID>
<name>N_in0</name></connection>
<connection>
<GID>163</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-79.5,98,-69</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<connection>
<GID>47</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>69,-98.5,69,-98.5</points>
<connection>
<GID>43</GID>
<name>A_greater_B</name></connection>
<connection>
<GID>165</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-102.5,69,-102.5</points>
<connection>
<GID>43</GID>
<name>A_less_B</name></connection>
<intersection>-102.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,-102.5,69,-102.5</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-100.5,69,-100.5</points>
<connection>
<GID>43</GID>
<name>A_equal_B</name></connection>
<intersection>-100.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,-100.5,69,-100.5</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-105.5,102.5,-99</points>
<intersection>-105.5 1</intersection>
<intersection>-99 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100.5,-105.5,102.5,-105.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>102.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>102.5,-99,104,-99</points>
<connection>
<GID>24</GID>
<name>carry_out</name></connection>
<intersection>102.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-96,133,-91</points>
<connection>
<GID>25</GID>
<name>IN_B_0</name></connection>
<intersection>-91 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>105,-91,105,-81.5</points>
<connection>
<GID>72</GID>
<name>N_in1</name></connection>
<intersection>-91 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>98,-91,133,-91</points>
<intersection>98 7</intersection>
<intersection>105 1</intersection>
<intersection>133 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>98,-96.5,98,-91</points>
<connection>
<GID>22</GID>
<name>IN_B_0</name></connection>
<intersection>-91 2</intersection></vsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-90.5,104,-81.5</points>
<connection>
<GID>71</GID>
<name>N_in1</name></connection>
<intersection>-90.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>132,-96,132,-90.5</points>
<connection>
<GID>25</GID>
<name>IN_B_1</name></connection>
<intersection>-90.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>97,-90.5,132,-90.5</points>
<intersection>97 7</intersection>
<intersection>104 0</intersection>
<intersection>132 1</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>97,-96.5,97,-90.5</points>
<connection>
<GID>22</GID>
<name>IN_B_1</name></connection>
<intersection>-90.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>131,-96,131,-90</points>
<connection>
<GID>25</GID>
<name>IN_B_2</name></connection>
<intersection>-90 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>103,-90,103,-81.5</points>
<connection>
<GID>53</GID>
<name>N_in1</name></connection>
<intersection>-90 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>96,-90,131,-90</points>
<intersection>96 7</intersection>
<intersection>103 1</intersection>
<intersection>131 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>96,-96.5,96,-90</points>
<connection>
<GID>22</GID>
<name>IN_B_2</name></connection>
<intersection>-90 2</intersection></vsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-89.5,102,-81.5</points>
<connection>
<GID>51</GID>
<name>N_in1</name></connection>
<intersection>-89.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>130,-96,130,-89.5</points>
<connection>
<GID>25</GID>
<name>IN_B_3</name></connection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>95,-89.5,130,-89.5</points>
<intersection>95 7</intersection>
<intersection>102 0</intersection>
<intersection>130 1</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>95,-96.5,95,-89.5</points>
<connection>
<GID>22</GID>
<name>IN_B_3</name></connection>
<intersection>-89.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117,-96,117,-89</points>
<connection>
<GID>24</GID>
<name>IN_B_0</name></connection>
<intersection>-89 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>101,-89,101,-81.5</points>
<connection>
<GID>50</GID>
<name>N_in1</name></connection>
<intersection>-89 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>82,-89,117,-89</points>
<intersection>82 7</intersection>
<intersection>101 1</intersection>
<intersection>117 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>82,-96.5,82,-89</points>
<connection>
<GID>43</GID>
<name>IN_B_0</name></connection>
<intersection>-89 2</intersection></vsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100,-88.5,100,-81.5</points>
<connection>
<GID>49</GID>
<name>N_in1</name></connection>
<intersection>-88.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>116,-96,116,-88.5</points>
<connection>
<GID>24</GID>
<name>IN_B_1</name></connection>
<intersection>-88.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>81,-88.5,116,-88.5</points>
<intersection>81 7</intersection>
<intersection>100 0</intersection>
<intersection>116 1</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>81,-96.5,81,-88.5</points>
<connection>
<GID>43</GID>
<name>IN_B_1</name></connection>
<intersection>-88.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-96,115,-88</points>
<connection>
<GID>24</GID>
<name>IN_B_2</name></connection>
<intersection>-88 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>99,-88,99,-81.5</points>
<connection>
<GID>48</GID>
<name>N_in1</name></connection>
<intersection>-88 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>80,-88,115,-88</points>
<intersection>80 7</intersection>
<intersection>99 1</intersection>
<intersection>115 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>80,-96.5,80,-88</points>
<connection>
<GID>43</GID>
<name>IN_B_2</name></connection>
<intersection>-88 2</intersection></vsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98,-87.5,98,-81.5</points>
<connection>
<GID>47</GID>
<name>N_in1</name></connection>
<intersection>-87.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>114,-96,114,-87.5</points>
<connection>
<GID>24</GID>
<name>IN_B_3</name></connection>
<intersection>-87.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>79,-87.5,114,-87.5</points>
<intersection>79 4</intersection>
<intersection>98 0</intersection>
<intersection>114 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>79,-96.5,79,-87.5</points>
<connection>
<GID>43</GID>
<name>IN_B_3</name></connection>
<intersection>-87.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-120,12,89.5</points>
<connection>
<GID>67</GID>
<name>N_in0</name></connection>
<connection>
<GID>59</GID>
<name>N_in1</name></connection>
<intersection>-81 10</intersection>
<intersection>-34.5 8</intersection>
<intersection>4 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>12,4,26,4</points>
<connection>
<GID>52</GID>
<name>IN_2</name></connection>
<intersection>12 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>12,-34.5,26,-34.5</points>
<connection>
<GID>121</GID>
<name>IN_2</name></connection>
<intersection>12 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>12,-81,48.5,-81</points>
<intersection>12 0</intersection>
<intersection>30.5 12</intersection>
<intersection>48.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>48.5,-81,48.5,-77.5</points>
<connection>
<GID>223</GID>
<name>IN_2</name></connection>
<intersection>-81 10</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>30.5,-81,30.5,-77.5</points>
<connection>
<GID>224</GID>
<name>IN_2</name></connection>
<intersection>-81 10</intersection></vsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-120,9,89.5</points>
<connection>
<GID>64</GID>
<name>N_in0</name></connection>
<connection>
<GID>56</GID>
<name>N_in1</name></connection>
<intersection>-79.5 9</intersection>
<intersection>-31.5 8</intersection>
<intersection>7 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>9,7,26,7</points>
<connection>
<GID>52</GID>
<name>IN_5</name></connection>
<intersection>9 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>9,-31.5,26,-31.5</points>
<connection>
<GID>121</GID>
<name>IN_5</name></connection>
<intersection>9 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>9,-79.5,45.5,-79.5</points>
<intersection>9 0</intersection>
<intersection>27.5 11</intersection>
<intersection>45.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>45.5,-79.5,45.5,-77.5</points>
<connection>
<GID>223</GID>
<name>IN_5</name></connection>
<intersection>-79.5 9</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>27.5,-79.5,27.5,-77.5</points>
<connection>
<GID>224</GID>
<name>IN_5</name></connection>
<intersection>-79.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-120,14,89.5</points>
<connection>
<GID>69</GID>
<name>N_in0</name></connection>
<connection>
<GID>61</GID>
<name>N_in1</name></connection>
<intersection>-82 10</intersection>
<intersection>-36.5 8</intersection>
<intersection>2 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>14,2,26,2</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>14,-36.5,26,-36.5</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>14,-82,50.5,-82</points>
<intersection>14 0</intersection>
<intersection>32.5 12</intersection>
<intersection>50.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>50.5,-82,50.5,-77.5</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>-82 10</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>32.5,-82,32.5,-77.5</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>-82 10</intersection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-120,10,89.5</points>
<connection>
<GID>65</GID>
<name>N_in0</name></connection>
<connection>
<GID>57</GID>
<name>N_in1</name></connection>
<intersection>-80 9</intersection>
<intersection>-32.5 8</intersection>
<intersection>6 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>10,6,26,6</points>
<connection>
<GID>52</GID>
<name>IN_4</name></connection>
<intersection>10 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>10,-32.5,26,-32.5</points>
<connection>
<GID>121</GID>
<name>IN_4</name></connection>
<intersection>10 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>10,-80,46.5,-80</points>
<intersection>10 0</intersection>
<intersection>28.5 11</intersection>
<intersection>46.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>46.5,-80,46.5,-77.5</points>
<connection>
<GID>223</GID>
<name>IN_4</name></connection>
<intersection>-80 9</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>28.5,-80,28.5,-77.5</points>
<connection>
<GID>224</GID>
<name>IN_4</name></connection>
<intersection>-80 9</intersection></vsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-120,11,89.5</points>
<connection>
<GID>66</GID>
<name>N_in0</name></connection>
<connection>
<GID>58</GID>
<name>N_in1</name></connection>
<intersection>-80.5 10</intersection>
<intersection>-33.5 8</intersection>
<intersection>5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>11,5,26,5</points>
<connection>
<GID>52</GID>
<name>IN_3</name></connection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>11,-33.5,26,-33.5</points>
<connection>
<GID>121</GID>
<name>IN_3</name></connection>
<intersection>11 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>11,-80.5,47.5,-80.5</points>
<intersection>11 0</intersection>
<intersection>29.5 12</intersection>
<intersection>47.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>47.5,-80.5,47.5,-77.5</points>
<connection>
<GID>223</GID>
<name>IN_3</name></connection>
<intersection>-80.5 10</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>29.5,-80.5,29.5,-77.5</points>
<connection>
<GID>224</GID>
<name>IN_3</name></connection>
<intersection>-80.5 10</intersection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-120,8,89.5</points>
<connection>
<GID>63</GID>
<name>N_in0</name></connection>
<connection>
<GID>55</GID>
<name>N_in1</name></connection>
<intersection>-79 9</intersection>
<intersection>-30.5 8</intersection>
<intersection>8 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>8,8,26,8</points>
<connection>
<GID>52</GID>
<name>IN_6</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>8,-30.5,26,-30.5</points>
<connection>
<GID>121</GID>
<name>IN_6</name></connection>
<intersection>8 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>8,-79,44.5,-79</points>
<intersection>8 0</intersection>
<intersection>26.5 11</intersection>
<intersection>44.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>44.5,-79,44.5,-77.5</points>
<connection>
<GID>223</GID>
<name>IN_6</name></connection>
<intersection>-79 9</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>26.5,-79,26.5,-77.5</points>
<connection>
<GID>224</GID>
<name>IN_6</name></connection>
<intersection>-79 9</intersection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-120,13,89.5</points>
<connection>
<GID>68</GID>
<name>N_in0</name></connection>
<connection>
<GID>60</GID>
<name>N_in1</name></connection>
<intersection>-81.5 9</intersection>
<intersection>-35.5 8</intersection>
<intersection>3 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>13,3,26,3</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>13,-35.5,26,-35.5</points>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>13,-81.5,49.5,-81.5</points>
<intersection>13 0</intersection>
<intersection>31.5 11</intersection>
<intersection>49.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>49.5,-81.5,49.5,-77.5</points>
<connection>
<GID>223</GID>
<name>IN_1</name></connection>
<intersection>-81.5 9</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>31.5,-81.5,31.5,-77.5</points>
<connection>
<GID>224</GID>
<name>IN_1</name></connection>
<intersection>-81.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,-120,7,89.5</points>
<connection>
<GID>62</GID>
<name>N_in0</name></connection>
<connection>
<GID>54</GID>
<name>N_in1</name></connection>
<intersection>-78.5 9</intersection>
<intersection>-29.5 8</intersection>
<intersection>9 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>7,9,26,9</points>
<connection>
<GID>52</GID>
<name>IN_7</name></connection>
<intersection>7 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>7,-29.5,26,-29.5</points>
<connection>
<GID>121</GID>
<name>IN_7</name></connection>
<intersection>7 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>7,-78.5,43.5,-78.5</points>
<intersection>7 0</intersection>
<intersection>25.5 11</intersection>
<intersection>43.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>43.5,-78.5,43.5,-77.5</points>
<connection>
<GID>223</GID>
<name>IN_7</name></connection>
<intersection>-78.5 9</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>25.5,-78.5,25.5,-77.5</points>
<connection>
<GID>224</GID>
<name>IN_7</name></connection>
<intersection>-78.5 9</intersection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,-96,126,-86</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-86 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>93,-86,93,-81.5</points>
<connection>
<GID>120</GID>
<name>N_in1</name></connection>
<intersection>-86 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>91,-86,126,-86</points>
<intersection>91 4</intersection>
<intersection>93 1</intersection>
<intersection>126 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>91,-96.5,91,-86</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-86 2</intersection></vsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,-85.5,92,-81.5</points>
<connection>
<GID>119</GID>
<name>N_in1</name></connection>
<intersection>-85.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>125,-96,125,-85.5</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>-85.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>90,-85.5,125,-85.5</points>
<intersection>90 4</intersection>
<intersection>92 0</intersection>
<intersection>125 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>90,-96.5,90,-85.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>-85.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,-96,124,-85</points>
<connection>
<GID>25</GID>
<name>IN_2</name></connection>
<intersection>-85 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>91,-85,91,-81.5</points>
<connection>
<GID>118</GID>
<name>N_in1</name></connection>
<intersection>-85 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>89,-85,124,-85</points>
<intersection>89 4</intersection>
<intersection>91 1</intersection>
<intersection>124 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>89,-96.5,89,-85</points>
<connection>
<GID>22</GID>
<name>IN_2</name></connection>
<intersection>-85 2</intersection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-84.5,90,-81.5</points>
<connection>
<GID>90</GID>
<name>N_in1</name></connection>
<intersection>-84.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>123,-96,123,-84.5</points>
<connection>
<GID>25</GID>
<name>IN_3</name></connection>
<intersection>-84.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>88,-84.5,123,-84.5</points>
<intersection>88 4</intersection>
<intersection>90 0</intersection>
<intersection>123 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>88,-96.5,88,-84.5</points>
<connection>
<GID>22</GID>
<name>IN_3</name></connection>
<intersection>-84.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-96,110,-84</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-84 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>89,-84,89,-81.5</points>
<connection>
<GID>84</GID>
<name>N_in1</name></connection>
<intersection>-84 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>75,-84,110,-84</points>
<intersection>75 4</intersection>
<intersection>89 1</intersection>
<intersection>110 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>75,-96.5,75,-84</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>-84 2</intersection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-83.5,88,-81.5</points>
<connection>
<GID>83</GID>
<name>N_in1</name></connection>
<intersection>-83.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>109,-96,109,-83.5</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>-83.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>74,-83.5,109,-83.5</points>
<intersection>74 4</intersection>
<intersection>88 0</intersection>
<intersection>109 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>74,-96.5,74,-83.5</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>-83.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-96,108,-83</points>
<connection>
<GID>24</GID>
<name>IN_2</name></connection>
<intersection>-83 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>87,-83,87,-81.5</points>
<connection>
<GID>75</GID>
<name>N_in1</name></connection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>73,-83,108,-83</points>
<intersection>73 4</intersection>
<intersection>87 1</intersection>
<intersection>108 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>73,-96.5,73,-83</points>
<connection>
<GID>43</GID>
<name>IN_2</name></connection>
<intersection>-83 2</intersection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-82.5,86,-81.5</points>
<connection>
<GID>73</GID>
<name>N_in1</name></connection>
<intersection>-82.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>107,-96,107,-82.5</points>
<connection>
<GID>24</GID>
<name>IN_3</name></connection>
<intersection>-82.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>72,-82.5,107,-82.5</points>
<intersection>72 4</intersection>
<intersection>86 0</intersection>
<intersection>107 1</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>72,-96.5,72,-82.5</points>
<connection>
<GID>43</GID>
<name>IN_3</name></connection>
<intersection>-82.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-99,136,-99</points>
<connection>
<GID>25</GID>
<name>carry_in</name></connection>
<connection>
<GID>169</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,11,29,12.5</points>
<connection>
<GID>52</GID>
<name>load</name></connection>
<intersection>12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,12.5,29,12.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-3.5,31,0</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<connection>
<GID>52</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103,-108,103,-101</points>
<intersection>-108 2</intersection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103,-101,104,-101</points>
<connection>
<GID>24</GID>
<name>overflow</name></connection>
<intersection>103 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>100.5,-108,103,-108</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>103 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,12,81.5,12</points>
<connection>
<GID>70</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>78</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,2,90,10</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,2,114,2</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>65.5 4</intersection>
<intersection>90 0</intersection>
<intersection>114 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>114,2,114,10</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>2 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>65.5,2,65.5,10</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>2 1</intersection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,3,89,10</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>3 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,3,113,3</points>
<connection>
<GID>52</GID>
<name>OUT_1</name></connection>
<intersection>64.5 4</intersection>
<intersection>89 0</intersection>
<intersection>113 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>113,3,113,10</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>3 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>64.5,3,64.5,10</points>
<connection>
<GID>81</GID>
<name>IN_1</name></connection>
<intersection>3 1</intersection></vsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,4,88,10</points>
<connection>
<GID>70</GID>
<name>IN_2</name></connection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,4,112,4</points>
<connection>
<GID>52</GID>
<name>OUT_2</name></connection>
<intersection>63.5 4</intersection>
<intersection>88 0</intersection>
<intersection>112 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>112,4,112,10</points>
<connection>
<GID>79</GID>
<name>IN_2</name></connection>
<intersection>4 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>63.5,4,63.5,10</points>
<connection>
<GID>81</GID>
<name>IN_2</name></connection>
<intersection>4 1</intersection></vsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,5,87,10</points>
<connection>
<GID>70</GID>
<name>IN_3</name></connection>
<intersection>5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,5,111,5</points>
<connection>
<GID>52</GID>
<name>OUT_3</name></connection>
<intersection>62.5 4</intersection>
<intersection>87 0</intersection>
<intersection>111 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>111,5,111,10</points>
<connection>
<GID>79</GID>
<name>IN_3</name></connection>
<intersection>5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>62.5,5,62.5,10</points>
<connection>
<GID>81</GID>
<name>IN_3</name></connection>
<intersection>5 1</intersection></vsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,6,86,10</points>
<connection>
<GID>70</GID>
<name>IN_4</name></connection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,6,110,6</points>
<connection>
<GID>52</GID>
<name>OUT_4</name></connection>
<intersection>61.5 4</intersection>
<intersection>86 0</intersection>
<intersection>110 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>110,6,110,10</points>
<connection>
<GID>79</GID>
<name>IN_4</name></connection>
<intersection>6 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>61.5,6,61.5,10</points>
<connection>
<GID>81</GID>
<name>IN_4</name></connection>
<intersection>6 1</intersection></vsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,7,85,10</points>
<connection>
<GID>70</GID>
<name>IN_5</name></connection>
<intersection>7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,7,109,7</points>
<connection>
<GID>52</GID>
<name>OUT_5</name></connection>
<intersection>60.5 4</intersection>
<intersection>85 0</intersection>
<intersection>109 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>109,7,109,10</points>
<connection>
<GID>79</GID>
<name>IN_5</name></connection>
<intersection>7 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>60.5,7,60.5,10</points>
<connection>
<GID>81</GID>
<name>IN_5</name></connection>
<intersection>7 1</intersection></vsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,8,84,10</points>
<connection>
<GID>70</GID>
<name>IN_6</name></connection>
<intersection>8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,8,108,8</points>
<connection>
<GID>52</GID>
<name>OUT_6</name></connection>
<intersection>59.5 5</intersection>
<intersection>84 0</intersection>
<intersection>108 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>108,8,108,10</points>
<connection>
<GID>79</GID>
<name>IN_6</name></connection>
<intersection>8 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>59.5,8,59.5,10</points>
<connection>
<GID>81</GID>
<name>IN_6</name></connection>
<intersection>8 1</intersection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,9,107,9</points>
<connection>
<GID>52</GID>
<name>OUT_7</name></connection>
<intersection>58.5 8</intersection>
<intersection>83 4</intersection>
<intersection>107 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>83,9,83,10</points>
<connection>
<GID>70</GID>
<name>IN_7</name></connection>
<intersection>9 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>107,9,107,10</points>
<connection>
<GID>79</GID>
<name>IN_7</name></connection>
<intersection>9 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>58.5,9,58.5,10</points>
<connection>
<GID>81</GID>
<name>IN_7</name></connection>
<intersection>9 1</intersection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,12,105.5,12</points>
<connection>
<GID>79</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>80</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,12,57,12</points>
<connection>
<GID>81</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>82</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,14,65.5,14</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<connection>
<GID>85</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,14,64.5,19</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<connection>
<GID>81</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,14,63.5,14</points>
<connection>
<GID>81</GID>
<name>OUT_2</name></connection>
<connection>
<GID>87</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,14,61.5,14</points>
<connection>
<GID>81</GID>
<name>OUT_4</name></connection>
<connection>
<GID>88</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,14,59.5,14</points>
<connection>
<GID>81</GID>
<name>OUT_6</name></connection>
<connection>
<GID>89</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>111,-116,115,-116</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>115 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>115,-116,115,-116</points>
<connection>
<GID>171</GID>
<name>ENABLE_0</name></connection>
<intersection>-116 1</intersection></vsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,14,58.5,19</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<connection>
<GID>81</GID>
<name>OUT_7</name></connection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,14,60.5,19</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<connection>
<GID>81</GID>
<name>OUT_5</name></connection></vsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,14,62.5,19</points>
<connection>
<GID>81</GID>
<name>OUT_3</name></connection>
<connection>
<GID>91</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,14,90,14</points>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<connection>
<GID>94</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,14,88,14</points>
<connection>
<GID>70</GID>
<name>OUT_2</name></connection>
<connection>
<GID>95</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,14,86,14</points>
<connection>
<GID>70</GID>
<name>OUT_4</name></connection>
<connection>
<GID>96</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,14,84,14</points>
<connection>
<GID>70</GID>
<name>OUT_6</name></connection>
<connection>
<GID>97</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,14,89,24.5</points>
<connection>
<GID>70</GID>
<name>OUT_1</name></connection>
<connection>
<GID>98</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,14,87,24.5</points>
<connection>
<GID>70</GID>
<name>OUT_3</name></connection>
<connection>
<GID>99</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-114,123.5,-114</points>
<connection>
<GID>171</GID>
<name>OUT_0</name></connection>
<connection>
<GID>173</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-114,122.5,-109</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<connection>
<GID>171</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,14,83,24.5</points>
<connection>
<GID>70</GID>
<name>OUT_7</name></connection>
<connection>
<GID>101</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,14,85,24.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<connection>
<GID>70</GID>
<name>OUT_5</name></connection></vsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,14,112,14</points>
<connection>
<GID>79</GID>
<name>OUT_2</name></connection>
<connection>
<GID>103</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,14,114,14</points>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection>
<connection>
<GID>102</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,14,110,14</points>
<connection>
<GID>79</GID>
<name>OUT_4</name></connection>
<connection>
<GID>104</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,14,108,14</points>
<connection>
<GID>79</GID>
<name>OUT_6</name></connection>
<connection>
<GID>105</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,91.5,12,91.5</points>
<connection>
<GID>59</GID>
<name>N_in0</name></connection>
<connection>
<GID>112</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,91.5,14,91.5</points>
<connection>
<GID>61</GID>
<name>N_in0</name></connection>
<connection>
<GID>110</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,91.5,10,91.5</points>
<connection>
<GID>57</GID>
<name>N_in0</name></connection>
<connection>
<GID>113</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,91.5,8,91.5</points>
<connection>
<GID>55</GID>
<name>N_in0</name></connection>
<connection>
<GID>114</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,91.5,13,96.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<connection>
<GID>60</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,91.5,11,96.5</points>
<connection>
<GID>58</GID>
<name>N_in0</name></connection>
<connection>
<GID>115</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,91.5,9,96.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<connection>
<GID>56</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7,91.5,7,96.5</points>
<connection>
<GID>54</GID>
<name>N_in0</name></connection>
<connection>
<GID>117</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-114,121.5,-114</points>
<connection>
<GID>171</GID>
<name>OUT_2</name></connection>
<connection>
<GID>175</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-27.5,29,-26</points>
<connection>
<GID>121</GID>
<name>load</name></connection>
<intersection>-26 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>28.5,-26,29,-26</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-41.5,31,-38.5</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<connection>
<GID>121</GID>
<name>clear</name></connection></vsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-26.5,81.5,-26.5</points>
<connection>
<GID>122</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>126</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-36.5,90,-28.5</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-36.5,114,-36.5</points>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection>
<intersection>65.5 4</intersection>
<intersection>90 0</intersection>
<intersection>114 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>114,-36.5,114,-28.5</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>-36.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>65.5,-36.5,65.5,-28.5</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<intersection>-36.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-35.5,89,-28.5</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-35.5,113,-35.5</points>
<connection>
<GID>121</GID>
<name>OUT_1</name></connection>
<intersection>64.5 4</intersection>
<intersection>89 0</intersection>
<intersection>113 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>113,-35.5,113,-28.5</points>
<connection>
<GID>127</GID>
<name>IN_1</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>64.5,-35.5,64.5,-28.5</points>
<connection>
<GID>129</GID>
<name>IN_1</name></connection>
<intersection>-35.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-34.5,88,-28.5</points>
<connection>
<GID>122</GID>
<name>IN_2</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-34.5,112,-34.5</points>
<connection>
<GID>121</GID>
<name>OUT_2</name></connection>
<intersection>63.5 4</intersection>
<intersection>88 0</intersection>
<intersection>112 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>112,-34.5,112,-28.5</points>
<connection>
<GID>127</GID>
<name>IN_2</name></connection>
<intersection>-34.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>63.5,-34.5,63.5,-28.5</points>
<connection>
<GID>129</GID>
<name>IN_2</name></connection>
<intersection>-34.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-33.5,87,-28.5</points>
<connection>
<GID>122</GID>
<name>IN_3</name></connection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-33.5,111,-33.5</points>
<connection>
<GID>121</GID>
<name>OUT_3</name></connection>
<intersection>62.5 4</intersection>
<intersection>87 0</intersection>
<intersection>111 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>111,-33.5,111,-28.5</points>
<connection>
<GID>127</GID>
<name>IN_3</name></connection>
<intersection>-33.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>62.5,-33.5,62.5,-28.5</points>
<connection>
<GID>129</GID>
<name>IN_3</name></connection>
<intersection>-33.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-32.5,86,-28.5</points>
<connection>
<GID>122</GID>
<name>IN_4</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-32.5,110,-32.5</points>
<connection>
<GID>121</GID>
<name>OUT_4</name></connection>
<intersection>61.5 4</intersection>
<intersection>86 0</intersection>
<intersection>110 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>110,-32.5,110,-28.5</points>
<connection>
<GID>127</GID>
<name>IN_4</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>61.5,-32.5,61.5,-28.5</points>
<connection>
<GID>129</GID>
<name>IN_4</name></connection>
<intersection>-32.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-31.5,85,-28.5</points>
<connection>
<GID>122</GID>
<name>IN_5</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-31.5,109,-31.5</points>
<connection>
<GID>121</GID>
<name>OUT_5</name></connection>
<intersection>60.5 4</intersection>
<intersection>85 0</intersection>
<intersection>109 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>109,-31.5,109,-28.5</points>
<connection>
<GID>127</GID>
<name>IN_5</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>60.5,-31.5,60.5,-28.5</points>
<connection>
<GID>129</GID>
<name>IN_5</name></connection>
<intersection>-31.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-30.5,84,-28.5</points>
<connection>
<GID>122</GID>
<name>IN_6</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-30.5,108,-30.5</points>
<connection>
<GID>121</GID>
<name>OUT_6</name></connection>
<intersection>59.5 5</intersection>
<intersection>84 0</intersection>
<intersection>108 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>108,-30.5,108,-28.5</points>
<connection>
<GID>127</GID>
<name>IN_6</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>59.5,-30.5,59.5,-28.5</points>
<connection>
<GID>129</GID>
<name>IN_6</name></connection>
<intersection>-30.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-29.5,107,-29.5</points>
<connection>
<GID>121</GID>
<name>OUT_7</name></connection>
<intersection>58.5 8</intersection>
<intersection>83 4</intersection>
<intersection>107 5</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>83,-29.5,83,-28.5</points>
<connection>
<GID>122</GID>
<name>IN_7</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>107,-29.5,107,-28.5</points>
<connection>
<GID>127</GID>
<name>IN_7</name></connection>
<intersection>-29.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>58.5,-29.5,58.5,-28.5</points>
<connection>
<GID>129</GID>
<name>IN_7</name></connection>
<intersection>-29.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105.5,-26.5,105.5,-26.5</points>
<connection>
<GID>127</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>128</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-26.5,57,-26.5</points>
<connection>
<GID>129</GID>
<name>ENABLE_0</name></connection>
<connection>
<GID>130</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-24.5,65.5,-24.5</points>
<connection>
<GID>129</GID>
<name>OUT_0</name></connection>
<connection>
<GID>131</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-24.5,64.5,-19.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<connection>
<GID>129</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-24.5,63.5,-24.5</points>
<connection>
<GID>129</GID>
<name>OUT_2</name></connection>
<connection>
<GID>133</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-24.5,61.5,-24.5</points>
<connection>
<GID>129</GID>
<name>OUT_4</name></connection>
<connection>
<GID>134</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-24.5,59.5,-24.5</points>
<connection>
<GID>129</GID>
<name>OUT_6</name></connection>
<connection>
<GID>135</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-24.5,58.5,-19.5</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<connection>
<GID>129</GID>
<name>OUT_7</name></connection></vsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-24.5,60.5,-19.5</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<connection>
<GID>129</GID>
<name>OUT_5</name></connection></vsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-24.5,62.5,-19.5</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<connection>
<GID>129</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-24.5,90,-24.5</points>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<connection>
<GID>139</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-24.5,88,-24.5</points>
<connection>
<GID>122</GID>
<name>OUT_2</name></connection>
<connection>
<GID>140</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-24.5,86,-24.5</points>
<connection>
<GID>122</GID>
<name>OUT_4</name></connection>
<connection>
<GID>141</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-24.5,84,-24.5</points>
<connection>
<GID>122</GID>
<name>OUT_6</name></connection>
<connection>
<GID>142</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-24.5,89,-14</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<connection>
<GID>122</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-24.5,87,-14</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<connection>
<GID>122</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-24.5,83,-14</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<connection>
<GID>122</GID>
<name>OUT_7</name></connection></vsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-24.5,85,-14</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<connection>
<GID>122</GID>
<name>OUT_5</name></connection></vsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-24.5,112,-24.5</points>
<connection>
<GID>127</GID>
<name>OUT_2</name></connection>
<connection>
<GID>148</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,-24.5,114,-24.5</points>
<connection>
<GID>127</GID>
<name>OUT_0</name></connection>
<connection>
<GID>147</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110,-24.5,110,-24.5</points>
<connection>
<GID>127</GID>
<name>OUT_4</name></connection>
<connection>
<GID>149</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>108,-24.5,108,-24.5</points>
<connection>
<GID>127</GID>
<name>OUT_6</name></connection>
<connection>
<GID>150</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-39.5,29,-38.5</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<connection>
<GID>121</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-1,29,0</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<connection>
<GID>52</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-7.5,-28,-7.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<connection>
<GID>159</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-114,119.5,-114</points>
<connection>
<GID>171</GID>
<name>OUT_4</name></connection>
<connection>
<GID>176</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-114,117.5,-114</points>
<connection>
<GID>171</GID>
<name>OUT_6</name></connection>
<connection>
<GID>177</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-114,116.5,-109</points>
<connection>
<GID>171</GID>
<name>OUT_7</name></connection>
<connection>
<GID>180</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-114,118.5,-109</points>
<connection>
<GID>171</GID>
<name>OUT_5</name></connection>
<connection>
<GID>179</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120.5,-114,120.5,-109</points>
<connection>
<GID>171</GID>
<name>OUT_3</name></connection>
<connection>
<GID>178</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-119,123.5,-118</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>-119 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>129.5,-119,129.5,-104</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>-119 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>123.5,-119,129.5,-119</points>
<intersection>123.5 0</intersection>
<intersection>129.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>164</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122.5,-119.5,122.5,-118</points>
<connection>
<GID>171</GID>
<name>IN_1</name></connection>
<intersection>-119.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>128.5,-119.5,128.5,-104</points>
<connection>
<GID>25</GID>
<name>OUT_1</name></connection>
<intersection>-119.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>122.5,-119.5,128.5,-119.5</points>
<intersection>122.5 0</intersection>
<intersection>128.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>165</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-120,121.5,-118</points>
<connection>
<GID>171</GID>
<name>IN_2</name></connection>
<intersection>-120 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>127.5,-120,127.5,-104</points>
<connection>
<GID>25</GID>
<name>OUT_2</name></connection>
<intersection>-120 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>121.5,-120,127.5,-120</points>
<intersection>121.5 0</intersection>
<intersection>127.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>166</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126.5,-120.5,126.5,-104</points>
<connection>
<GID>25</GID>
<name>OUT_3</name></connection>
<intersection>-120.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>120.5,-120.5,120.5,-118</points>
<connection>
<GID>171</GID>
<name>IN_3</name></connection>
<intersection>-120.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>120.5,-120.5,126.5,-120.5</points>
<intersection>120.5 1</intersection>
<intersection>126.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>167</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-120.5,119.5,-118</points>
<connection>
<GID>171</GID>
<name>IN_4</name></connection>
<intersection>-120.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>113.5,-120.5,113.5,-104</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>-120.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>113.5,-120.5,119.5,-120.5</points>
<intersection>113.5 1</intersection>
<intersection>119.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>168</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-120,112.5,-104</points>
<connection>
<GID>24</GID>
<name>OUT_1</name></connection>
<intersection>-120 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>118.5,-120,118.5,-118</points>
<connection>
<GID>171</GID>
<name>IN_5</name></connection>
<intersection>-120 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>112.5,-120,118.5,-120</points>
<intersection>112.5 0</intersection>
<intersection>118.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>169</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117.5,-119.5,117.5,-118</points>
<connection>
<GID>171</GID>
<name>IN_6</name></connection>
<intersection>-119.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>111.5,-119.5,111.5,-104</points>
<connection>
<GID>24</GID>
<name>OUT_2</name></connection>
<intersection>-119.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>111.5,-119.5,117.5,-119.5</points>
<intersection>111.5 1</intersection>
<intersection>117.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>170</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-119,110.5,-104</points>
<connection>
<GID>24</GID>
<name>OUT_3</name></connection>
<intersection>-119 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>116.5,-119,116.5,-118</points>
<connection>
<GID>171</GID>
<name>IN_7</name></connection>
<intersection>-119 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>110.5,-119,116.5,-119</points>
<intersection>110.5 0</intersection>
<intersection>116.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>179</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>26.5,-71.5,26.5,-71.5</points>
<connection>
<GID>209</GID>
<name>N_in0</name></connection>
<connection>
<GID>193</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>180</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>28.5,-71.5,28.5,-71.5</points>
<connection>
<GID>211</GID>
<name>N_in0</name></connection>
<connection>
<GID>192</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>181</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30.5,-71.5,30.5,-71.5</points>
<connection>
<GID>213</GID>
<name>N_in0</name></connection>
<connection>
<GID>191</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>182</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>32.5,-71.5,32.5,-71.5</points>
<connection>
<GID>215</GID>
<name>N_in0</name></connection>
<connection>
<GID>190</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>183</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-71.5,31.5,-61</points>
<connection>
<GID>214</GID>
<name>N_in0</name></connection>
<connection>
<GID>194</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>184</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-71.5,29.5,-61</points>
<connection>
<GID>212</GID>
<name>N_in0</name></connection>
<connection>
<GID>195</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>185</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-71.5,27.5,-61</points>
<connection>
<GID>210</GID>
<name>N_in0</name></connection>
<connection>
<GID>196</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>186</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-71.5,25.5,-61</points>
<connection>
<GID>208</GID>
<name>N_in0</name></connection>
<connection>
<GID>197</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>187</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>44.5,-71.5,44.5,-71.5</points>
<connection>
<GID>201</GID>
<name>N_in0</name></connection>
<connection>
<GID>217</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>188</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>46.5,-71.5,46.5,-71.5</points>
<connection>
<GID>203</GID>
<name>N_in0</name></connection>
<connection>
<GID>216</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>189</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>48.5,-71.5,48.5,-71.5</points>
<connection>
<GID>205</GID>
<name>N_in0</name></connection>
<connection>
<GID>199</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>190</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>50.5,-71.5,50.5,-71.5</points>
<connection>
<GID>207</GID>
<name>N_in0</name></connection>
<connection>
<GID>198</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>191</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-71.5,49.5,-61</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<connection>
<GID>206</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>192</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47.5,-71.5,47.5,-61</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<connection>
<GID>204</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>193</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-71.5,45.5,-61</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<connection>
<GID>202</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>194</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-71.5,43.5,-61</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<connection>
<GID>200</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>195</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>50.5,-73.5,50.5,-73.5</points>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection>
<connection>
<GID>207</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>196</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>43.5,-73.5,43.5,-73.5</points>
<connection>
<GID>223</GID>
<name>OUT_7</name></connection>
<connection>
<GID>200</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>197</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>44.5,-73.5,44.5,-73.5</points>
<connection>
<GID>223</GID>
<name>OUT_6</name></connection>
<connection>
<GID>201</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>198</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>47.5,-73.5,47.5,-73.5</points>
<connection>
<GID>223</GID>
<name>OUT_3</name></connection>
<connection>
<GID>204</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>199</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>49.5,-73.5,49.5,-73.5</points>
<connection>
<GID>223</GID>
<name>OUT_1</name></connection>
<connection>
<GID>206</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>200</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>45.5,-73.5,45.5,-73.5</points>
<connection>
<GID>223</GID>
<name>OUT_5</name></connection>
<connection>
<GID>202</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>201</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>46.5,-73.5,46.5,-73.5</points>
<connection>
<GID>223</GID>
<name>OUT_4</name></connection>
<connection>
<GID>203</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>202</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>48.5,-73.5,48.5,-73.5</points>
<connection>
<GID>223</GID>
<name>OUT_2</name></connection>
<connection>
<GID>205</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>203</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>25.5,-73.5,25.5,-73.5</points>
<connection>
<GID>224</GID>
<name>OUT_7</name></connection>
<connection>
<GID>208</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>204</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>27.5,-73.5,27.5,-73.5</points>
<connection>
<GID>224</GID>
<name>OUT_5</name></connection>
<connection>
<GID>210</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>205</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>28.5,-73.5,28.5,-73.5</points>
<connection>
<GID>224</GID>
<name>OUT_4</name></connection>
<connection>
<GID>211</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>206</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>29.5,-73.5,29.5,-73.5</points>
<connection>
<GID>224</GID>
<name>OUT_3</name></connection>
<connection>
<GID>212</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>207</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>30.5,-73.5,30.5,-73.5</points>
<connection>
<GID>224</GID>
<name>OUT_2</name></connection>
<connection>
<GID>213</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>208</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>32.5,-73.5,32.5,-73.5</points>
<connection>
<GID>224</GID>
<name>OUT_0</name></connection>
<connection>
<GID>215</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>209</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>31.5,-73.5,31.5,-73.5</points>
<connection>
<GID>224</GID>
<name>OUT_1</name></connection>
<connection>
<GID>214</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>210</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>26.5,-73.5,26.5,-73.5</points>
<connection>
<GID>224</GID>
<name>OUT_6</name></connection>
<connection>
<GID>209</GID>
<name>N_in1</name></connection></hsegment></shape></wire>
<wire>
<ID>211</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-75.5,41,-74.5</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41,-75.5,42,-75.5</points>
<connection>
<GID>223</GID>
<name>ENABLE_0</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>212</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-75.5,23,-74.5</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<intersection>-75.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-75.5,24,-75.5</points>
<connection>
<GID>224</GID>
<name>ENABLE_0</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>218</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43.5,-121.5,-43.5,-70.5</points>
<intersection>-121.5 6</intersection>
<intersection>-104.5 7</intersection>
<intersection>-87.5 4</intersection>
<intersection>-73.5 2</intersection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-43.5,-70.5,-36,-70.5</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>-43.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-52,-73.5,-43.5,-73.5</points>
<connection>
<GID>241</GID>
<name>OUT_0</name></connection>
<intersection>-43.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-43.5,-87.5,-36,-87.5</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>-43.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-43.5,-121.5,-36,-121.5</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>-43.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-43.5,-104.5,-36,-104.5</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>-43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>219</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44,-120.5,-44,-69.5</points>
<intersection>-120.5 8</intersection>
<intersection>-103.5 6</intersection>
<intersection>-86.5 4</intersection>
<intersection>-71.5 1</intersection>
<intersection>-69.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-52,-71.5,-44,-71.5</points>
<connection>
<GID>241</GID>
<name>OUT_1</name></connection>
<intersection>-44 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-44,-69.5,-36,-69.5</points>
<connection>
<GID>234</GID>
<name>IN_1</name></connection>
<intersection>-44 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-44,-86.5,-36,-86.5</points>
<connection>
<GID>235</GID>
<name>IN_1</name></connection>
<intersection>-44 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-44,-103.5,-36,-103.5</points>
<connection>
<GID>247</GID>
<name>IN_1</name></connection>
<intersection>-44 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-44,-120.5,-36,-120.5</points>
<connection>
<GID>248</GID>
<name>IN_1</name></connection>
<intersection>-44 0</intersection></hsegment></shape></wire>
<wire>
<ID>220</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-44.5,-119.5,-44.5,-68.5</points>
<intersection>-119.5 8</intersection>
<intersection>-102.5 6</intersection>
<intersection>-85.5 4</intersection>
<intersection>-69.5 2</intersection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-44.5,-68.5,-36,-68.5</points>
<connection>
<GID>234</GID>
<name>IN_2</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-52,-69.5,-44.5,-69.5</points>
<connection>
<GID>241</GID>
<name>OUT_2</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-44.5,-85.5,-36,-85.5</points>
<connection>
<GID>235</GID>
<name>IN_2</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-44.5,-102.5,-36,-102.5</points>
<connection>
<GID>247</GID>
<name>IN_2</name></connection>
<intersection>-44.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>-44.5,-119.5,-36,-119.5</points>
<connection>
<GID>248</GID>
<name>IN_2</name></connection>
<intersection>-44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>221</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-45,-118.5,-45,-67.5</points>
<intersection>-118.5 9</intersection>
<intersection>-101.5 7</intersection>
<intersection>-84.5 4</intersection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-52,-67.5,-36,-67.5</points>
<connection>
<GID>234</GID>
<name>IN_3</name></connection>
<connection>
<GID>241</GID>
<name>OUT_3</name></connection>
<intersection>-45 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-45,-84.5,-36,-84.5</points>
<connection>
<GID>235</GID>
<name>IN_3</name></connection>
<intersection>-45 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-45,-101.5,-36,-101.5</points>
<connection>
<GID>247</GID>
<name>IN_3</name></connection>
<intersection>-45 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-45,-118.5,-36,-118.5</points>
<connection>
<GID>248</GID>
<name>IN_3</name></connection>
<intersection>-45 0</intersection></hsegment></shape></wire>
<wire>
<ID>224</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63.5,-85.5,-63.5,-73.5</points>
<intersection>-85.5 2</intersection>
<intersection>-73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64,-73.5,-63.5,-73.5</points>
<connection>
<GID>242</GID>
<name>OUT_0</name></connection>
<intersection>-63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-63.5,-85.5,-61.5,-85.5</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>-63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>225</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,-84.5,-63,-71.5</points>
<intersection>-84.5 2</intersection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64,-71.5,-63,-71.5</points>
<connection>
<GID>242</GID>
<name>OUT_1</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-63,-84.5,-61.5,-84.5</points>
<connection>
<GID>244</GID>
<name>IN_1</name></connection>
<intersection>-63 0</intersection></hsegment></shape></wire>
<wire>
<ID>226</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62,-82.5,-62,-82</points>
<connection>
<GID>246</GID>
<name>OUT_0</name></connection>
<intersection>-82.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-62,-82.5,-61.5,-82.5</points>
<connection>
<GID>244</GID>
<name>ENABLE</name></connection>
<intersection>-62 0</intersection></hsegment></shape></wire>
<wire>
<ID>227</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,-106.5,-46,-85.5</points>
<intersection>-106.5 1</intersection>
<intersection>-85.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-46,-106.5,-36,-106.5</points>
<connection>
<GID>248</GID>
<name>ENABLE</name></connection>
<intersection>-46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-55.5,-85.5,-46,-85.5</points>
<connection>
<GID>244</GID>
<name>OUT_0</name></connection>
<intersection>-46 0</intersection></hsegment></shape></wire>
<wire>
<ID>228</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-45.5,-89.5,-45.5,-84.5</points>
<intersection>-89.5 1</intersection>
<intersection>-84.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,-89.5,-36,-89.5</points>
<connection>
<GID>247</GID>
<name>ENABLE</name></connection>
<intersection>-45.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-55.5,-84.5,-45.5,-84.5</points>
<connection>
<GID>244</GID>
<name>OUT_1</name></connection>
<intersection>-45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>229</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-45.5,-83.5,-45.5,-72.5</points>
<intersection>-83.5 2</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,-72.5,-36,-72.5</points>
<connection>
<GID>235</GID>
<name>ENABLE</name></connection>
<intersection>-45.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-55.5,-83.5,-45.5,-83.5</points>
<connection>
<GID>244</GID>
<name>OUT_2</name></connection>
<intersection>-45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>230</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-46,-82.5,-46,-55.5</points>
<intersection>-82.5 2</intersection>
<intersection>-55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-46,-55.5,-36,-55.5</points>
<connection>
<GID>234</GID>
<name>ENABLE</name></connection>
<intersection>-46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-55.5,-82.5,-46,-82.5</points>
<connection>
<GID>244</GID>
<name>OUT_3</name></connection>
<intersection>-46 0</intersection></hsegment></shape></wire>
<wire>
<ID>236</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-30,-103.5,-16,-103.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<connection>
<GID>247</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>237</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-87.5,-30,-87.5</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<connection>
<GID>235</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>239</ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-30,-55.5,-30,-55.5</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<connection>
<GID>234</GID>
<name>OUT_15</name></connection></hsegment></shape></wire>
<wire>
<ID>240</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-104.5,-30,-104.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<connection>
<GID>247</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>241</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195.5,-121,195.5,-70</points>
<intersection>-121 6</intersection>
<intersection>-104 7</intersection>
<intersection>-87 4</intersection>
<intersection>-73 2</intersection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>195.5,-70,203,-70</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>187,-73,195.5,-73</points>
<connection>
<GID>256</GID>
<name>OUT_0</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>195.5,-87,203,-87</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>195.5,-121,203,-121</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<intersection>195.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>195.5,-104,203,-104</points>
<connection>
<GID>260</GID>
<name>IN_0</name></connection>
<intersection>195.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>242</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>195,-120,195,-69</points>
<intersection>-120 8</intersection>
<intersection>-103 6</intersection>
<intersection>-86 4</intersection>
<intersection>-71 1</intersection>
<intersection>-69 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>187,-71,195,-71</points>
<connection>
<GID>256</GID>
<name>OUT_1</name></connection>
<intersection>195 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>195,-69,203,-69</points>
<connection>
<GID>254</GID>
<name>IN_1</name></connection>
<intersection>195 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>195,-86,203,-86</points>
<connection>
<GID>255</GID>
<name>IN_1</name></connection>
<intersection>195 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>195,-103,203,-103</points>
<connection>
<GID>260</GID>
<name>IN_1</name></connection>
<intersection>195 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>195,-120,203,-120</points>
<connection>
<GID>261</GID>
<name>IN_1</name></connection>
<intersection>195 0</intersection></hsegment></shape></wire>
<wire>
<ID>243</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194.5,-119,194.5,-68</points>
<intersection>-119 8</intersection>
<intersection>-102 6</intersection>
<intersection>-85 4</intersection>
<intersection>-69 2</intersection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>194.5,-68,203,-68</points>
<connection>
<GID>254</GID>
<name>IN_2</name></connection>
<intersection>194.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>187,-69,194.5,-69</points>
<connection>
<GID>256</GID>
<name>OUT_2</name></connection>
<intersection>194.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>194.5,-85,203,-85</points>
<connection>
<GID>255</GID>
<name>IN_2</name></connection>
<intersection>194.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>194.5,-102,203,-102</points>
<connection>
<GID>260</GID>
<name>IN_2</name></connection>
<intersection>194.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>194.5,-119,203,-119</points>
<connection>
<GID>261</GID>
<name>IN_2</name></connection>
<intersection>194.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>244</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>194,-118,194,-67</points>
<intersection>-118 9</intersection>
<intersection>-101 7</intersection>
<intersection>-84 4</intersection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>187,-67,203,-67</points>
<connection>
<GID>254</GID>
<name>IN_3</name></connection>
<connection>
<GID>256</GID>
<name>OUT_3</name></connection>
<intersection>194 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>194,-84,203,-84</points>
<connection>
<GID>255</GID>
<name>IN_3</name></connection>
<intersection>194 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>194,-101,203,-101</points>
<connection>
<GID>260</GID>
<name>IN_3</name></connection>
<intersection>194 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>194,-118,203,-118</points>
<connection>
<GID>261</GID>
<name>IN_3</name></connection>
<intersection>194 0</intersection></hsegment></shape></wire>
<wire>
<ID>245</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175.5,-85,175.5,-73</points>
<intersection>-85 2</intersection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175,-73,175.5,-73</points>
<connection>
<GID>257</GID>
<name>OUT_0</name></connection>
<intersection>175.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>175.5,-85,177.5,-85</points>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>175.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>246</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>176,-84,176,-71</points>
<intersection>-84 2</intersection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175,-71,176,-71</points>
<connection>
<GID>257</GID>
<name>OUT_1</name></connection>
<intersection>176 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>176,-84,177.5,-84</points>
<connection>
<GID>258</GID>
<name>IN_1</name></connection>
<intersection>176 0</intersection></hsegment></shape></wire>
<wire>
<ID>247</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>177,-82,177,-81.5</points>
<connection>
<GID>259</GID>
<name>OUT_0</name></connection>
<intersection>-82 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>177,-82,177.5,-82</points>
<connection>
<GID>258</GID>
<name>ENABLE</name></connection>
<intersection>177 0</intersection></hsegment></shape></wire>
<wire>
<ID>248</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193,-106,193,-85</points>
<intersection>-106 1</intersection>
<intersection>-85 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>193,-106,203,-106</points>
<connection>
<GID>261</GID>
<name>ENABLE</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>183.5,-85,193,-85</points>
<connection>
<GID>258</GID>
<name>OUT_0</name></connection>
<intersection>193 0</intersection></hsegment></shape></wire>
<wire>
<ID>249</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193.5,-89,193.5,-84</points>
<intersection>-89 1</intersection>
<intersection>-84 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>193.5,-89,203,-89</points>
<connection>
<GID>260</GID>
<name>ENABLE</name></connection>
<intersection>193.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>183.5,-84,193.5,-84</points>
<connection>
<GID>258</GID>
<name>OUT_1</name></connection>
<intersection>193.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>250</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193.5,-83,193.5,-72</points>
<intersection>-83 2</intersection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>193.5,-72,203,-72</points>
<connection>
<GID>255</GID>
<name>ENABLE</name></connection>
<intersection>193.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>183.5,-83,193.5,-83</points>
<connection>
<GID>258</GID>
<name>OUT_2</name></connection>
<intersection>193.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>251</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193,-82,193,-55</points>
<intersection>-82 2</intersection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>193,-55,203,-55</points>
<connection>
<GID>254</GID>
<name>ENABLE</name></connection>
<intersection>193 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>183.5,-82,193,-82</points>
<connection>
<GID>258</GID>
<name>OUT_3</name></connection>
<intersection>193 0</intersection></hsegment></shape></wire>
<wire>
<ID>252</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264,-120,264,-69</points>
<intersection>-120 6</intersection>
<intersection>-103 7</intersection>
<intersection>-86 4</intersection>
<intersection>-72 2</intersection>
<intersection>-69 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>264,-69,271.5,-69</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<intersection>264 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>255.5,-72,264,-72</points>
<connection>
<GID>264</GID>
<name>OUT_0</name></connection>
<intersection>264 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>264,-86,271.5,-86</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<intersection>264 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>264,-120,271.5,-120</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>264 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>264,-103,271.5,-103</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<intersection>264 0</intersection></hsegment></shape></wire>
<wire>
<ID>253</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>263.5,-119,263.5,-68</points>
<intersection>-119 8</intersection>
<intersection>-102 6</intersection>
<intersection>-85 4</intersection>
<intersection>-70 1</intersection>
<intersection>-68 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255.5,-70,263.5,-70</points>
<connection>
<GID>264</GID>
<name>OUT_1</name></connection>
<intersection>263.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>263.5,-68,271.5,-68</points>
<connection>
<GID>262</GID>
<name>IN_1</name></connection>
<intersection>263.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>263.5,-85,271.5,-85</points>
<connection>
<GID>263</GID>
<name>IN_1</name></connection>
<intersection>263.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>263.5,-102,271.5,-102</points>
<connection>
<GID>268</GID>
<name>IN_1</name></connection>
<intersection>263.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>263.5,-119,271.5,-119</points>
<connection>
<GID>269</GID>
<name>IN_1</name></connection>
<intersection>263.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>254</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>263,-118,263,-67</points>
<intersection>-118 8</intersection>
<intersection>-101 6</intersection>
<intersection>-84 4</intersection>
<intersection>-68 2</intersection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>263,-67,271.5,-67</points>
<connection>
<GID>262</GID>
<name>IN_2</name></connection>
<intersection>263 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>255.5,-68,263,-68</points>
<connection>
<GID>264</GID>
<name>OUT_2</name></connection>
<intersection>263 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>263,-84,271.5,-84</points>
<connection>
<GID>263</GID>
<name>IN_2</name></connection>
<intersection>263 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>263,-101,271.5,-101</points>
<connection>
<GID>268</GID>
<name>IN_2</name></connection>
<intersection>263 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>263,-118,271.5,-118</points>
<connection>
<GID>269</GID>
<name>IN_2</name></connection>
<intersection>263 0</intersection></hsegment></shape></wire>
<wire>
<ID>255</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262.5,-117,262.5,-66</points>
<intersection>-117 9</intersection>
<intersection>-100 7</intersection>
<intersection>-83 4</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>255.5,-66,271.5,-66</points>
<connection>
<GID>262</GID>
<name>IN_3</name></connection>
<connection>
<GID>264</GID>
<name>OUT_3</name></connection>
<intersection>262.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>262.5,-83,271.5,-83</points>
<connection>
<GID>263</GID>
<name>IN_3</name></connection>
<intersection>262.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>262.5,-100,271.5,-100</points>
<connection>
<GID>268</GID>
<name>IN_3</name></connection>
<intersection>262.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>262.5,-117,271.5,-117</points>
<connection>
<GID>269</GID>
<name>IN_3</name></connection>
<intersection>262.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>256</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244,-84,244,-72</points>
<intersection>-84 2</intersection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>243.5,-72,244,-72</points>
<connection>
<GID>265</GID>
<name>OUT_0</name></connection>
<intersection>244 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>244,-84,246,-84</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<intersection>244 0</intersection></hsegment></shape></wire>
<wire>
<ID>257</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>244.5,-83,244.5,-70</points>
<intersection>-83 2</intersection>
<intersection>-70 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>243.5,-70,244.5,-70</points>
<connection>
<GID>265</GID>
<name>OUT_1</name></connection>
<intersection>244.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>244.5,-83,246,-83</points>
<connection>
<GID>266</GID>
<name>IN_1</name></connection>
<intersection>244.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>258</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>245.5,-81,245.5,-80.5</points>
<connection>
<GID>267</GID>
<name>OUT_0</name></connection>
<intersection>-81 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>245.5,-81,246,-81</points>
<connection>
<GID>266</GID>
<name>ENABLE</name></connection>
<intersection>245.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>259</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261.5,-105,261.5,-84</points>
<intersection>-105 1</intersection>
<intersection>-84 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261.5,-105,271.5,-105</points>
<connection>
<GID>269</GID>
<name>ENABLE</name></connection>
<intersection>261.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>252,-84,261.5,-84</points>
<connection>
<GID>266</GID>
<name>OUT_0</name></connection>
<intersection>261.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>260</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262,-88,262,-83</points>
<intersection>-88 1</intersection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>262,-88,271.5,-88</points>
<connection>
<GID>268</GID>
<name>ENABLE</name></connection>
<intersection>262 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>252,-83,262,-83</points>
<connection>
<GID>266</GID>
<name>OUT_1</name></connection>
<intersection>262 0</intersection></hsegment></shape></wire>
<wire>
<ID>261</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>262,-82,262,-71</points>
<intersection>-82 2</intersection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>262,-71,271.5,-71</points>
<connection>
<GID>263</GID>
<name>ENABLE</name></connection>
<intersection>262 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>252,-82,262,-82</points>
<connection>
<GID>266</GID>
<name>OUT_2</name></connection>
<intersection>262 0</intersection></hsegment></shape></wire>
<wire>
<ID>262</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>261.5,-81,261.5,-54</points>
<intersection>-81 2</intersection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>261.5,-54,271.5,-54</points>
<connection>
<GID>262</GID>
<name>ENABLE</name></connection>
<intersection>261.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>252,-81,261.5,-81</points>
<connection>
<GID>266</GID>
<name>OUT_3</name></connection>
<intersection>261.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>263</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>209,-104,209,-104</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<connection>
<GID>260</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>264</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>209,-103,224,-103</points>
<connection>
<GID>260</GID>
<name>OUT_1</name></connection>
<connection>
<GID>271</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>265</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277.5,-103,277.5,-103</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<connection>
<GID>268</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>266</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>277.5,-102,292,-102</points>
<connection>
<GID>268</GID>
<name>OUT_1</name></connection>
<connection>
<GID>273</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>267</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>277.5,-69,277.5,-69</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<connection>
<GID>262</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>268</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>209,-70,209,-70</points>
<connection>
<GID>254</GID>
<name>OUT_0</name></connection>
<connection>
<GID>275</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>269</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-70.5,-30,-70.5</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<connection>
<GID>234</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>270</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-74.5,-26.5,-74.5,-26.5</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<connection>
<GID>278</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>272</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-74.5,-24.5,-74.5,-24.5</points>
<connection>
<GID>277</GID>
<name>IN_2</name></connection>
<connection>
<GID>280</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>273</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-74.5,-22.5,-74.5,-22.5</points>
<connection>
<GID>277</GID>
<name>IN_4</name></connection>
<connection>
<GID>281</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>274</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-74.5,-20.5,-74.5,-20.5</points>
<connection>
<GID>277</GID>
<name>IN_6</name></connection>
<connection>
<GID>282</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>275</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80,-19.5,-74.5,-19.5</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<connection>
<GID>277</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>276</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80,-21.5,-74.5,-21.5</points>
<connection>
<GID>277</GID>
<name>IN_5</name></connection>
<connection>
<GID>284</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>277</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80,-23.5,-74.5,-23.5</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<connection>
<GID>277</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>278</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80,-25.5,-74.5,-25.5</points>
<connection>
<GID>277</GID>
<name>IN_1</name></connection>
<connection>
<GID>279</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>279</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-24.5,-28,-24.5</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<connection>
<GID>287</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>280</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-29,-28,-29</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<connection>
<GID>290</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>281</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-32,-28,-32</points>
<connection>
<GID>291</GID>
<name>OUT_0</name></connection>
<connection>
<GID>289</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>282</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-24.5,107,-14</points>
<connection>
<GID>127</GID>
<name>OUT_7</name></connection>
<connection>
<GID>154</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>283</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,-24.5,109,-14</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<connection>
<GID>127</GID>
<name>OUT_5</name></connection></vsegment></shape></wire>
<wire>
<ID>284</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-24.5,111,-14</points>
<connection>
<GID>127</GID>
<name>OUT_3</name></connection>
<connection>
<GID>152</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>285</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,-24.5,113,-14</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<connection>
<GID>127</GID>
<name>OUT_1</name></connection></vsegment></shape></wire>
<wire>
<ID>286</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,14,107,24.5</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<connection>
<GID>79</GID>
<name>OUT_7</name></connection></vsegment></shape></wire>
<wire>
<ID>287</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>109,14,109,24.5</points>
<connection>
<GID>79</GID>
<name>OUT_5</name></connection>
<connection>
<GID>108</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>288</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,14,111,24.5</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<connection>
<GID>79</GID>
<name>OUT_3</name></connection></vsegment></shape></wire>
<wire>
<ID>289</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>113,14,113,24.5</points>
<connection>
<GID>79</GID>
<name>OUT_1</name></connection>
<connection>
<GID>106</GID>
<name>IN_0</name></connection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-8.42641e-006,43.329,594.646,-288.687</PageViewport></page 1>
<page 2>
<PageViewport>-8.42641e-006,43.329,594.646,-288.687</PageViewport></page 2>
<page 3>
<PageViewport>-8.42641e-006,43.329,594.646,-288.687</PageViewport></page 3>
<page 4>
<PageViewport>-8.42641e-006,43.329,594.646,-288.687</PageViewport></page 4>
<page 5>
<PageViewport>-8.42641e-006,43.329,594.646,-288.687</PageViewport></page 5>
<page 6>
<PageViewport>-8.42641e-006,43.329,594.646,-288.687</PageViewport></page 6>
<page 7>
<PageViewport>-8.42641e-006,43.329,594.646,-288.687</PageViewport></page 7>
<page 8>
<PageViewport>-8.42641e-006,43.329,594.646,-288.687</PageViewport></page 8>
<page 9>
<PageViewport>-8.42641e-006,43.329,594.646,-288.687</PageViewport></page 9></circuit>